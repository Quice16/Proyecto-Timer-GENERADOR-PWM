VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO timer_pwm_interface
  CLASS BLOCK ;
  FOREIGN timer_pwm_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 94.445 BY 105.165 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.020 10.640 16.620 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.380 89.020 21.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.720 10.640 13.320 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.080 89.020 18.680 ;
    END
  END VPWR
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 101.165 55.110 105.165 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 64.640 94.445 65.240 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 101.165 67.990 105.165 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 101.165 61.550 105.165 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 68.040 94.445 68.640 ;
    END
  END addr[4]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END clk
  PIN irq_timer
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 64.490 101.165 64.770 105.165 ;
    END
  END irq_timer
  PIN outa
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END outa
  PIN outb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END outb
  PIN rdata[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 90.445 78.240 94.445 78.840 ;
    END
  END rdata[0]
  PIN rdata[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 90.445 61.240 94.445 61.840 ;
    END
  END rdata[1]
  PIN rdata[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 90.445 57.840 94.445 58.440 ;
    END
  END rdata[2]
  PIN rdata[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 58.050 101.165 58.330 105.165 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 38.730 101.165 39.010 105.165 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 41.950 101.165 42.230 105.165 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 35.510 101.165 35.790 105.165 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 45.170 101.165 45.450 105.165 ;
    END
  END rdata[7]
  PIN read_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 101.165 48.670 105.165 ;
    END
  END read_en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 90.445 17.040 94.445 17.640 ;
    END
  END rst
  PIN wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 71.440 94.445 72.040 ;
    END
  END wdata[0]
  PIN wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 54.440 94.445 55.040 ;
    END
  END wdata[1]
  PIN wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 47.640 94.445 48.240 ;
    END
  END wdata[2]
  PIN wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 90.445 51.040 94.445 51.640 ;
    END
  END wdata[3]
  PIN wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 101.165 29.350 105.165 ;
    END
  END wdata[4]
  PIN wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wdata[5]
  PIN wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wdata[6]
  PIN wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wdata[7]
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 101.165 51.890 105.165 ;
    END
  END write_en
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 88.970 92.565 ;
      LAYER li1 ;
        RECT 5.520 10.795 88.780 92.565 ;
      LAYER met1 ;
        RECT 4.210 10.640 88.780 92.720 ;
      LAYER met2 ;
        RECT 4.230 100.885 28.790 101.730 ;
        RECT 29.630 100.885 35.230 101.730 ;
        RECT 36.070 100.885 38.450 101.730 ;
        RECT 39.290 100.885 41.670 101.730 ;
        RECT 42.510 100.885 44.890 101.730 ;
        RECT 45.730 100.885 48.110 101.730 ;
        RECT 48.950 100.885 51.330 101.730 ;
        RECT 52.170 100.885 54.550 101.730 ;
        RECT 55.390 100.885 57.770 101.730 ;
        RECT 58.610 100.885 60.990 101.730 ;
        RECT 61.830 100.885 64.210 101.730 ;
        RECT 65.050 100.885 67.430 101.730 ;
        RECT 68.270 100.885 87.310 101.730 ;
        RECT 4.230 10.695 87.310 100.885 ;
      LAYER met3 ;
        RECT 3.990 86.040 90.445 92.645 ;
        RECT 4.400 84.640 90.445 86.040 ;
        RECT 3.990 79.240 90.445 84.640 ;
        RECT 3.990 77.840 90.045 79.240 ;
        RECT 3.990 75.840 90.445 77.840 ;
        RECT 4.400 74.440 90.445 75.840 ;
        RECT 3.990 72.440 90.445 74.440 ;
        RECT 3.990 71.040 90.045 72.440 ;
        RECT 3.990 69.040 90.445 71.040 ;
        RECT 3.990 67.640 90.045 69.040 ;
        RECT 3.990 65.640 90.445 67.640 ;
        RECT 4.400 64.240 90.045 65.640 ;
        RECT 3.990 62.240 90.445 64.240 ;
        RECT 3.990 60.840 90.045 62.240 ;
        RECT 3.990 58.840 90.445 60.840 ;
        RECT 3.990 57.440 90.045 58.840 ;
        RECT 3.990 55.440 90.445 57.440 ;
        RECT 4.400 54.040 90.045 55.440 ;
        RECT 3.990 52.040 90.445 54.040 ;
        RECT 3.990 50.640 90.045 52.040 ;
        RECT 3.990 48.640 90.445 50.640 ;
        RECT 3.990 47.240 90.045 48.640 ;
        RECT 3.990 41.840 90.445 47.240 ;
        RECT 4.400 40.440 90.445 41.840 ;
        RECT 3.990 38.440 90.445 40.440 ;
        RECT 4.400 37.040 90.445 38.440 ;
        RECT 3.990 18.040 90.445 37.040 ;
        RECT 3.990 16.640 90.045 18.040 ;
        RECT 3.990 10.715 90.445 16.640 ;
      LAYER met4 ;
        RECT 74.815 48.455 75.145 62.385 ;
  END
END timer_pwm_interface
END LIBRARY

