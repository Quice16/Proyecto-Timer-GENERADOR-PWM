* NGSPICE file created from timer_pwm_interface.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt timer_pwm_interface VGND VPWR addr[0] addr[1] addr[2] addr[3] addr[4] clk
+ irq_timer outa outb rdata[0] rdata[1] rdata[2] rdata[3] rdata[4] rdata[5] rdata[6]
+ rdata[7] read_en rst wdata[0] wdata[1] wdata[2] wdata[3] wdata[4] wdata[5] wdata[6]
+ wdata[7] write_en
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_294_ period\[7\] cnt\[7\] net2 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__mux2_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_363_ clknet_2_2__leaf_clk _057_ _032_ VGND VGND VPWR VPWR period\[3\] sky130_fd_sc_hd__dfrtp_1
X_346_ net7 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
XFILLER_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_277_ duty\[5\] _068_ _069_ duty\[4\] VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__o22a_1
XFILLER_5_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_200_ net14 period\[6\] _079_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__mux2_1
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_329_ net7 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR rdata[0] sky130_fd_sc_hd__buf_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_293_ _017_ net6 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nand2_2
X_362_ clknet_2_2__leaf_clk _056_ _031_ VGND VGND VPWR VPWR period\[2\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_12_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_345_ net7 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
X_276_ duty\[5\] _068_ _139_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ net7 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_259_ _113_ _106_ _093_ enable _125_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__o2111a_1
XFILLER_9_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR rdata[1] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_2_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_292_ _017_ net6 VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and2_2
XFILLER_26_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ clknet_2_2__leaf_clk _055_ _030_ VGND VGND VPWR VPWR period\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_344_ net7 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
X_275_ duty\[7\] _066_ _136_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ net15 duty\[7\] _077_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__mux2_1
X_327_ net7 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
X_258_ _068_ _123_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__xor2_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput22 net22 VGND VGND VPWR VPWR rdata[2] sky130_fd_sc_hd__buf_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ _017_ _074_ _152_ _115_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__o22ai_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_360_ clknet_2_3__leaf_clk _054_ _029_ VGND VGND VPWR VPWR period\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_343_ net7 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
X_274_ cnt\[5\] duty\[5\] VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ net16 _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand2_4
X_257_ _064_ _094_ _124_ _114_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nor4b_1
X_326_ net7 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ period\[2\] cnt\[2\] net2 VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__mux2_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput23 net23 VGND VGND VPWR VPWR rdata[3] sky130_fd_sc_hd__buf_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_290_ _017_ enable VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342_ net7 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
X_273_ duty\[7\] cnt\[7\] VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_187_ net1 _075_ _073_ net2 VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and4b_4
X_256_ _121_ _123_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ net7 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__bufinv_16
X_308_ net23 _153_ _164_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__o21a_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_239_ _108_ _109_ _089_ _091_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__o211ai_1
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput24 net24 VGND VGND VPWR VPWR rdata[4] sky130_fd_sc_hd__buf_1
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_341_ net7 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ cnt\[6\] duty\[6\] VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__nand2b_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_186_ net4 net5 VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_255_ _118_ _122_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__nand2_1
X_324_ net7 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_307_ _163_ _078_ _076_ duty\[3\] _154_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__a221o_1
X_238_ period\[5\] _068_ _108_ _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o22a_1
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VGND VPWR VPWR rdata[5] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_340_ net7 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__inv_2
X_271_ _132_ _133_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__a21o_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_323_ net7 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
X_185_ irq_timer_next VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__inv_2
X_254_ cnt\[4\] cnt\[3\] VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_28_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_306_ period\[3\] cnt\[3\] net2 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__mux2_1
X_237_ period\[4\] cnt\[4\] VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__and2_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput26 net26 VGND VGND VPWR VPWR rdata[6] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ _065_ cnt\[3\] _070_ duty\[2\] VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_322_ net7 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
X_184_ net7 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
X_253_ cnt\[3\] cnt\[2\] cnt\[1\] cnt\[0\] cnt\[4\] VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__a41o_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ net24 _153_ _162_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__o21a_1
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_236_ period\[4\] cnt\[4\] VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nor2_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_219_ _068_ period\[5\] VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__nand2_1
Xoutput27 net27 VGND VGND VPWR VPWR rdata[7] sky130_fd_sc_hd__buf_1
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_183_ net3 VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_252_ _113_ _106_ _093_ enable _120_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__o2111a_1
X_321_ net7 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
X_304_ _161_ _078_ _076_ duty\[4\] _154_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__a221o_1
X_235_ _104_ _098_ _105_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_218_ period\[4\] _069_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__o21ai_1
Xoutput17 net17 VGND VGND VPWR VPWR irq_timer sky130_fd_sc_hd__buf_1
XFILLER_7_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_320_ net20 _153_ _171_ _173_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__a2bb2oi_1
X_182_ cnt\[0\] VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ cnt\[3\] _118_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__xor2_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_303_ period\[4\] cnt\[4\] net2 VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__mux2_1
X_234_ _104_ _098_ _105_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_217_ period\[5\] cnt\[5\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand2b_1
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR outa sky130_fd_sc_hd__buf_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_181_ cnt\[1\] VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__inv_2
X_250_ _113_ _106_ _093_ enable _119_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__o2111a_1
X_379_ clknet_2_1__leaf_clk _047_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
X_302_ net25 _153_ _160_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__o21a_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ period\[2\] _070_ _099_ _101_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__o31a_1
XFILLER_29_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_216_ _082_ _083_ _086_ _087_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__nand4_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput19 net19 VGND VGND VPWR VPWR outb sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_17_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ cnt\[2\] VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__inv_2
X_378_ clknet_2_1__leaf_clk _046_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_301_ _159_ _078_ _076_ duty\[5\] _154_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__a221o_1
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_232_ _100_ _101_ _102_ _103_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_23_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_215_ cnt\[6\] period\[6\] VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_377_ clknet_2_0__leaf_clk _045_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
XFILLER_1_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ period\[5\] cnt\[5\] net2 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__mux2_1
X_231_ cnt\[2\] period\[2\] VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__nand2b_1
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_214_ cnt\[7\] period\[7\] VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ clknet_2_3__leaf_clk _044_ VGND VGND VPWR VPWR irq_timer_next sky130_fd_sc_hd__dfxtp_1
X_230_ period\[2\] cnt\[2\] VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__nand2b_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_359_ clknet_2_0__leaf_clk _007_ _028_ VGND VGND VPWR VPWR cnt\[7\] sky130_fd_sc_hd__dfrtp_2
Xinput2 addr[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_213_ _066_ period\[7\] VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__and2_1
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_375_ clknet_2_1__leaf_clk _043_ _016_ VGND VGND VPWR VPWR duty\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_358_ clknet_2_0__leaf_clk _006_ _027_ VGND VGND VPWR VPWR cnt\[6\] sky130_fd_sc_hd__dfrtp_4
Xinput3 addr[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ _142_ _149_ _148_ enable VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__o211a_1
XFILLER_19_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_212_ period\[7\] _066_ _067_ period\[6\] VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_27_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_374_ clknet_2_1__leaf_clk _042_ _015_ VGND VGND VPWR VPWR duty\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 addr[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_357_ clknet_2_0__leaf_clk _005_ _026_ VGND VGND VPWR VPWR cnt\[5\] sky130_fd_sc_hd__dfrtp_4
X_288_ _148_ _151_ _064_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_211_ period\[7\] cnt\[7\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_2_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_373_ clknet_2_1__leaf_clk _041_ _014_ VGND VGND VPWR VPWR duty\[5\] sky130_fd_sc_hd__dfstp_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 addr[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_287_ _138_ _141_ _147_ _150_ _137_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__o311a_1
X_356_ clknet_2_2__leaf_clk _004_ _025_ VGND VGND VPWR VPWR cnt\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_210_ period\[6\] cnt\[6\] VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2b_1
X_339_ net7 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__inv_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_372_ clknet_2_1__leaf_clk _040_ _013_ VGND VGND VPWR VPWR duty\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_286_ _066_ duty\[7\] duty\[6\] _067_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__a211o_1
X_355_ clknet_2_2__leaf_clk _003_ _024_ VGND VGND VPWR VPWR cnt\[3\] sky130_fd_sc_hd__dfrtp_4
Xinput6 read_en VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net7 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
X_269_ _071_ duty\[1\] duty\[2\] _070_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a22oi_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ clknet_2_3__leaf_clk _039_ _012_ VGND VGND VPWR VPWR duty\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_285_ _138_ _139_ _141_ _144_ _137_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__o311a_1
XFILLER_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_354_ clknet_2_2__leaf_clk _002_ _023_ VGND VGND VPWR VPWR cnt\[2\] sky130_fd_sc_hd__dfrtp_2
Xinput7 rst VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_12
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_337_ net7 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__inv_2
X_268_ duty\[1\] _071_ _072_ duty\[0\] VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o211ai_1
X_199_ net15 period\[7\] _079_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 wdata[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_13_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_370_ clknet_2_2__leaf_clk _038_ _011_ VGND VGND VPWR VPWR duty\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_284_ _135_ _140_ _141_ _146_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__nand4_1
X_353_ clknet_2_2__leaf_clk _001_ _022_ VGND VGND VPWR VPWR cnt\[1\] sky130_fd_sc_hd__dfrtp_4
Xinput8 wdata[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_336_ net7 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
X_198_ net2 net16 _078_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__nand3b_4
X_267_ _113_ _106_ _093_ enable _131_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__o2111a_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_319_ duty\[0\] _076_ _169_ _172_ _154_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_16_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 wdata[3] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_283_ _136_ _137_ _143_ _144_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__nand4_1
Xinput9 wdata[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_352_ clknet_2_2__leaf_clk _000_ _021_ VGND VGND VPWR VPWR cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_197_ net1 _075_ _073_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__and3_4
XFILLER_18_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ _129_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__nor2_1
X_335_ net7 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 wdata[4] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_318_ net2 net1 net4 net5 VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_249_ _117_ _118_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__nor2_1
XFILLER_20_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_351_ clknet_2_3__leaf_clk irq_timer_next _020_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_282_ cnt\[3\] _065_ _144_ _143_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__o2111a_1
XFILLER_14_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_334_ net7 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
X_196_ net8 duty\[0\] _077_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_265_ cnt\[6\] cnt\[5\] _118_ _122_ cnt\[7\] VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__a41oi_1
XTAP_TAPCELL_ROW_11_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_317_ _078_ _170_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__nand2_1
Xinput13 wdata[5] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_179_ cnt\[4\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__inv_2
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_248_ cnt\[2\] cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_281_ _069_ duty\[4\] VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__nand2_1
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ clknet_2_0__leaf_clk _009_ _019_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_195_ net9 duty\[1\] _077_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__mux2_1
X_333_ net7 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_264_ _066_ _127_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_316_ period\[0\] cnt\[0\] net2 VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__mux2_1
Xinput14 wdata[6] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_247_ cnt\[1\] cnt\[0\] cnt\[2\] VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_22_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_178_ cnt\[5\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__inv_2
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_280_ duty\[6\] cnt\[6\] VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__nand2b_1
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ net10 duty\[2\] _077_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__mux2_1
X_332_ net7 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
X_263_ _113_ _106_ _093_ enable _128_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_315_ enable net17 net3 VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__mux2_1
Xinput15 wdata[7] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_177_ cnt\[6\] VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__inv_2
X_246_ _113_ _106_ _093_ enable _116_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__o2111a_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_229_ period\[3\] cnt\[3\] VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nand2b_1
XFILLER_17_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ net11 duty\[3\] _077_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
X_331_ net7 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_262_ _126_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 write_en VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_314_ net21 _153_ _168_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__o21a_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_176_ cnt\[7\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__inv_2
X_245_ cnt\[1\] cnt\[0\] VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_228_ cnt\[3\] period\[3\] VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nand2b_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_192_ net12 duty\[4\] _077_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__mux2_1
XFILLER_25_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_330_ net7 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
X_261_ cnt\[6\] cnt\[5\] _118_ _122_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__nand4_1
XFILLER_11_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_313_ _167_ _078_ _076_ duty\[1\] _154_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__a221o_1
X_175_ duty\[3\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__inv_2
X_244_ _113_ _106_ _072_ enable _093_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__o2111a_1
XFILLER_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ cnt\[3\] period\[3\] VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__and2b_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_260_ cnt\[5\] _118_ _122_ cnt\[6\] VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a31o_1
X_191_ net13 duty\[5\] _077_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__mux2_1
XFILLER_17_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_312_ period\[1\] cnt\[1\] net2 VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__mux2_1
X_243_ _107_ _112_ _094_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__a21oi_1
X_174_ enable VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__inv_2
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_226_ _096_ _097_ _095_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_12_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_209_ enable net8 _081_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ net14 duty\[6\] _077_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__mux2_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ net22 _153_ _166_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__o21a_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_242_ _107_ _112_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__nand2_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_225_ cnt\[1\] period\[1\] VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__nand2b_1
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_208_ net16 _075_ _080_ _073_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__and4_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_310_ _165_ _078_ _076_ duty\[2\] _154_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__a221o_1
XFILLER_11_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ _088_ _091_ _110_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__nand3b_4
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_224_ cnt\[0\] period\[0\] VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nand2b_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_207_ net2 net1 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nor2_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_240_ _088_ _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__nor2_1
X_369_ clknet_2_3__leaf_clk _063_ _010_ VGND VGND VPWR VPWR duty\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_22_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_223_ period\[1\] cnt\[1\] VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__and2b_1
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_206_ net8 period\[0\] _079_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_299_ net26 _153_ _158_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__o21a_1
X_368_ clknet_2_3__leaf_clk _062_ _037_ VGND VGND VPWR VPWR duty\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_222_ _084_ _085_ _088_ _092_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__o22ai_1
X_205_ net9 period\[1\] _079_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__mux2_1
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_384_ clknet_2_3__leaf_clk _052_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ _157_ _078_ _076_ duty\[6\] _154_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__a221o_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_367_ clknet_2_0__leaf_clk _061_ _036_ VGND VGND VPWR VPWR period\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_221_ _084_ _085_ _088_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__o22a_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_204_ net10 period\[2\] _079_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__mux2_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_383_ clknet_2_3__leaf_clk _051_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_297_ period\[6\] cnt\[6\] net2 VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__mux2_1
X_366_ clknet_2_1__leaf_clk _060_ _035_ VGND VGND VPWR VPWR period\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ _090_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand2_1
X_349_ clknet_2_0__leaf_clk _008_ _018_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_23_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_203_ net11 period\[3\] _079_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_382_ clknet_2_3__leaf_clk _050_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_365_ clknet_2_1__leaf_clk _059_ _034_ VGND VGND VPWR VPWR period\[5\] sky130_fd_sc_hd__dfstp_1
XFILLER_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_296_ net27 _153_ _156_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__o21a_1
XFILLER_13_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ clknet_2_3__leaf_clk _053_ _017_ VGND VGND VPWR VPWR enable sky130_fd_sc_hd__dfrtp_4
X_279_ _066_ duty\[7\] VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_202_ net12 period\[4\] _079_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__mux2_1
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_381_ clknet_2_3__leaf_clk _049_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_364_ clknet_2_1__leaf_clk _058_ _033_ VGND VGND VPWR VPWR period\[4\] sky130_fd_sc_hd__dfrtp_1
X_295_ _155_ _078_ _076_ duty\[7\] _154_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__a221o_1
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_347_ net7 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
X_278_ _066_ duty\[7\] VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__and2_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_201_ net13 period\[5\] _079_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__mux2_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_380_ clknet_2_1__leaf_clk _048_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

