magic
tech sky130A
magscale 1 2
timestamp 1748585426
<< viali >>
rect 7205 18377 7239 18411
rect 7849 18377 7883 18411
rect 8493 18377 8527 18411
rect 9137 18377 9171 18411
rect 11713 18377 11747 18411
rect 13001 18377 13035 18411
rect 10517 18309 10551 18343
rect 2329 18241 2363 18275
rect 6101 18241 6135 18275
rect 6561 18241 6595 18275
rect 6837 18241 6871 18275
rect 7389 18241 7423 18275
rect 8033 18241 8067 18275
rect 8677 18241 8711 18275
rect 9321 18241 9355 18275
rect 9965 18241 9999 18275
rect 11069 18241 11103 18275
rect 11897 18241 11931 18275
rect 12357 18241 12391 18275
rect 13185 18241 13219 18275
rect 13645 18241 13679 18275
rect 10701 18105 10735 18139
rect 2421 18037 2455 18071
rect 5917 18037 5951 18071
rect 6377 18037 6411 18071
rect 6745 18037 6779 18071
rect 9781 18037 9815 18071
rect 11253 18037 11287 18071
rect 12541 18037 12575 18071
rect 13829 18037 13863 18071
rect 7113 17833 7147 17867
rect 12081 17833 12115 17867
rect 13921 17833 13955 17867
rect 1409 17697 1443 17731
rect 3801 17697 3835 17731
rect 14657 17697 14691 17731
rect 1777 17629 1811 17663
rect 4169 17629 4203 17663
rect 5733 17629 5767 17663
rect 7389 17629 7423 17663
rect 9229 17629 9263 17663
rect 10701 17629 10735 17663
rect 12173 17629 12207 17663
rect 14289 17629 14323 17663
rect 6000 17561 6034 17595
rect 7656 17561 7690 17595
rect 9496 17561 9530 17595
rect 10968 17561 11002 17595
rect 12449 17561 12483 17595
rect 14197 17561 14231 17595
rect 14924 17561 14958 17595
rect 3203 17493 3237 17527
rect 5595 17493 5629 17527
rect 8769 17493 8803 17527
rect 10609 17493 10643 17527
rect 16037 17493 16071 17527
rect 2053 17289 2087 17323
rect 2513 17289 2547 17323
rect 3985 17289 4019 17323
rect 4169 17289 4203 17323
rect 4537 17289 4571 17323
rect 4629 17289 4663 17323
rect 7757 17289 7791 17323
rect 7849 17289 7883 17323
rect 11529 17289 11563 17323
rect 13737 17289 13771 17323
rect 2421 17153 2455 17187
rect 3893 17153 3927 17187
rect 6377 17153 6411 17187
rect 6644 17153 6678 17187
rect 8033 17153 8067 17187
rect 8309 17153 8343 17187
rect 9321 17153 9355 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 10609 17153 10643 17187
rect 11713 17153 11747 17187
rect 11989 17153 12023 17187
rect 13369 17153 13403 17187
rect 13829 17153 13863 17187
rect 16313 17153 16347 17187
rect 17049 17153 17083 17187
rect 2697 17085 2731 17119
rect 4721 17085 4755 17119
rect 8217 17085 8251 17119
rect 9505 17085 9539 17119
rect 10517 17085 10551 17119
rect 13645 17085 13679 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 9413 17017 9447 17051
rect 9689 17017 9723 17051
rect 9873 17017 9907 17051
rect 9505 16949 9539 16983
rect 11897 16949 11931 16983
rect 13277 16949 13311 16983
rect 14197 16949 14231 16983
rect 16405 16949 16439 16983
rect 16681 16949 16715 16983
rect 6561 16745 6595 16779
rect 6929 16745 6963 16779
rect 9413 16745 9447 16779
rect 7021 16609 7055 16643
rect 9781 16609 9815 16643
rect 15669 16609 15703 16643
rect 15945 16609 15979 16643
rect 6745 16541 6779 16575
rect 9597 16541 9631 16575
rect 17417 16405 17451 16439
rect 14013 16201 14047 16235
rect 14841 16201 14875 16235
rect 14933 16201 14967 16235
rect 14105 16133 14139 16167
rect 2789 16065 2823 16099
rect 9505 16065 9539 16099
rect 9689 16065 9723 16099
rect 13829 16065 13863 16099
rect 13921 16065 13955 16099
rect 14197 16065 14231 16099
rect 14289 16065 14323 16099
rect 15117 16065 15151 16099
rect 15301 16065 15335 16099
rect 17233 16065 17267 16099
rect 9413 15997 9447 16031
rect 14749 15997 14783 16031
rect 2697 15861 2731 15895
rect 17417 15861 17451 15895
rect 3387 15657 3421 15691
rect 6929 15657 6963 15691
rect 7665 15657 7699 15691
rect 13645 15657 13679 15691
rect 13829 15657 13863 15691
rect 3801 15521 3835 15555
rect 8217 15521 8251 15555
rect 8309 15521 8343 15555
rect 11069 15521 11103 15555
rect 12173 15521 12207 15555
rect 12541 15521 12575 15555
rect 15945 15521 15979 15555
rect 1593 15453 1627 15487
rect 1961 15453 1995 15487
rect 5825 15453 5859 15487
rect 6285 15453 6319 15487
rect 6433 15453 6467 15487
rect 6769 15453 6803 15487
rect 7021 15453 7055 15487
rect 7114 15453 7148 15487
rect 7527 15453 7561 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13185 15453 13219 15487
rect 13553 15453 13587 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 4077 15385 4111 15419
rect 5733 15385 5767 15419
rect 6561 15385 6595 15419
rect 6653 15385 6687 15419
rect 7297 15385 7331 15419
rect 7389 15385 7423 15419
rect 9045 15385 9079 15419
rect 10793 15385 10827 15419
rect 11989 15385 12023 15419
rect 12633 15385 12667 15419
rect 13461 15385 13495 15419
rect 13829 15385 13863 15419
rect 16190 15385 16224 15419
rect 5549 15317 5583 15351
rect 7757 15317 7791 15351
rect 8125 15317 8159 15351
rect 11437 15317 11471 15351
rect 11621 15317 11655 15351
rect 12081 15317 12115 15351
rect 14197 15317 14231 15351
rect 17325 15317 17359 15351
rect 2237 15113 2271 15147
rect 2697 15113 2731 15147
rect 4537 15113 4571 15147
rect 4997 15113 5031 15147
rect 6929 15113 6963 15147
rect 9505 15113 9539 15147
rect 11897 15113 11931 15147
rect 12173 15113 12207 15147
rect 14565 15113 14599 15147
rect 15853 15113 15887 15147
rect 11621 15045 11655 15079
rect 11989 15045 12023 15079
rect 13001 15045 13035 15079
rect 1409 14977 1443 15011
rect 2605 14977 2639 15011
rect 4905 14977 4939 15011
rect 7297 14977 7331 15011
rect 7389 14977 7423 15011
rect 9597 14977 9631 15011
rect 10057 14977 10091 15011
rect 10701 14977 10735 15011
rect 11161 14977 11195 15011
rect 11805 14977 11839 15011
rect 12909 14977 12943 15011
rect 14381 14977 14415 15011
rect 14565 14977 14599 15011
rect 16037 14977 16071 15011
rect 2881 14909 2915 14943
rect 5181 14909 5215 14943
rect 7481 14909 7515 14943
rect 10977 14909 11011 14943
rect 12449 14909 12483 14943
rect 13185 14909 13219 14943
rect 16221 14909 16255 14943
rect 16313 14909 16347 14943
rect 1593 14841 1627 14875
rect 6653 14569 6687 14603
rect 17233 14569 17267 14603
rect 2329 14365 2363 14399
rect 4261 14365 4295 14399
rect 6009 14365 6043 14399
rect 6102 14365 6136 14399
rect 6285 14365 6319 14399
rect 6515 14365 6549 14399
rect 10701 14365 10735 14399
rect 10977 14365 11011 14399
rect 11345 14365 11379 14399
rect 17417 14365 17451 14399
rect 6377 14297 6411 14331
rect 2421 14229 2455 14263
rect 4353 14229 4387 14263
rect 6377 14025 6411 14059
rect 9045 14025 9079 14059
rect 11253 14025 11287 14059
rect 12541 14025 12575 14059
rect 14381 14025 14415 14059
rect 15117 14025 15151 14059
rect 17233 14025 17267 14059
rect 10885 13957 10919 13991
rect 3341 13889 3375 13923
rect 5135 13889 5169 13923
rect 6745 13889 6779 13923
rect 7932 13889 7966 13923
rect 9965 13889 9999 13923
rect 10609 13889 10643 13923
rect 10757 13889 10791 13923
rect 10977 13889 11011 13923
rect 11115 13889 11149 13923
rect 12633 13889 12667 13923
rect 14013 13889 14047 13923
rect 14473 13889 14507 13923
rect 14621 13889 14655 13923
rect 14749 13889 14783 13923
rect 14841 13889 14875 13923
rect 14938 13889 14972 13923
rect 15945 13889 15979 13923
rect 16129 13889 16163 13923
rect 17417 13889 17451 13923
rect 1409 13821 1443 13855
rect 1685 13821 1719 13855
rect 3157 13821 3191 13855
rect 3709 13821 3743 13855
rect 6837 13821 6871 13855
rect 6929 13821 6963 13855
rect 7665 13821 7699 13855
rect 10057 13821 10091 13855
rect 12817 13821 12851 13855
rect 13737 13821 13771 13855
rect 13921 13821 13955 13855
rect 16221 13821 16255 13855
rect 12173 13685 12207 13719
rect 15761 13685 15795 13719
rect 2145 13481 2179 13515
rect 3801 13481 3835 13515
rect 7941 13481 7975 13515
rect 8309 13481 8343 13515
rect 13277 13481 13311 13515
rect 14933 13481 14967 13515
rect 17233 13481 17267 13515
rect 2697 13345 2731 13379
rect 4445 13345 4479 13379
rect 8401 13345 8435 13379
rect 9045 13345 9079 13379
rect 11529 13345 11563 13379
rect 15853 13345 15887 13379
rect 1409 13277 1443 13311
rect 5641 13277 5675 13311
rect 8125 13277 8159 13311
rect 14289 13277 14323 13311
rect 14437 13277 14471 13311
rect 14565 13277 14599 13311
rect 14795 13277 14829 13311
rect 16109 13277 16143 13311
rect 2513 13209 2547 13243
rect 4169 13209 4203 13243
rect 4261 13209 4295 13243
rect 7389 13209 7423 13243
rect 9321 13209 9355 13243
rect 11805 13209 11839 13243
rect 14657 13209 14691 13243
rect 1593 13141 1627 13175
rect 2605 13141 2639 13175
rect 10793 13141 10827 13175
rect 7021 12937 7055 12971
rect 10057 12937 10091 12971
rect 13277 12937 13311 12971
rect 5733 12869 5767 12903
rect 6653 12869 6687 12903
rect 6745 12869 6779 12903
rect 4261 12801 4295 12835
rect 4353 12801 4387 12835
rect 4537 12801 4571 12835
rect 4629 12801 4663 12835
rect 6377 12801 6411 12835
rect 6470 12801 6504 12835
rect 6861 12801 6895 12835
rect 10425 12801 10459 12835
rect 10517 12801 10551 12835
rect 11805 12801 11839 12835
rect 13859 12801 13893 12835
rect 14013 12801 14047 12835
rect 14473 12801 14507 12835
rect 16681 12801 16715 12835
rect 17417 12801 17451 12835
rect 10701 12733 10735 12767
rect 17141 12733 17175 12767
rect 13645 12665 13679 12699
rect 4077 12597 4111 12631
rect 14565 12597 14599 12631
rect 16865 12597 16899 12631
rect 3157 12393 3191 12427
rect 7757 12393 7791 12427
rect 12541 12393 12575 12427
rect 4629 12325 4663 12359
rect 6561 12325 6595 12359
rect 7941 12325 7975 12359
rect 1409 12257 1443 12291
rect 6469 12257 6503 12291
rect 16681 12257 16715 12291
rect 3525 12189 3559 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 4813 12189 4847 12223
rect 4997 12189 5031 12223
rect 5548 12189 5582 12223
rect 5641 12189 5675 12223
rect 6008 12189 6042 12223
rect 6101 12189 6135 12223
rect 6929 12189 6963 12223
rect 7481 12189 7515 12223
rect 7573 12189 7607 12223
rect 7831 12189 7865 12223
rect 8125 12189 8159 12223
rect 8217 12189 8251 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 10701 12189 10735 12223
rect 12449 12189 12483 12223
rect 15577 12189 15611 12223
rect 15945 12189 15979 12223
rect 16865 12189 16899 12223
rect 1685 12121 1719 12155
rect 3433 12121 3467 12155
rect 7941 12121 7975 12155
rect 4353 12053 4387 12087
rect 5273 12053 5307 12087
rect 5733 12053 5767 12087
rect 7297 12053 7331 12087
rect 8401 12053 8435 12087
rect 10609 12053 10643 12087
rect 14151 12053 14185 12087
rect 16037 12053 16071 12087
rect 16405 12053 16439 12087
rect 16497 12053 16531 12087
rect 16957 12053 16991 12087
rect 2145 11849 2179 11883
rect 2605 11849 2639 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 7757 11849 7791 11883
rect 7849 11849 7883 11883
rect 12541 11849 12575 11883
rect 13093 11849 13127 11883
rect 14473 11849 14507 11883
rect 2513 11781 2547 11815
rect 8125 11781 8159 11815
rect 12173 11781 12207 11815
rect 14933 11781 14967 11815
rect 4261 11713 4295 11747
rect 4537 11713 4571 11747
rect 4721 11713 4755 11747
rect 5089 11713 5123 11747
rect 5181 11713 5215 11747
rect 5825 11713 5859 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 7665 11713 7699 11747
rect 8033 11713 8067 11747
rect 8401 11713 8435 11747
rect 8493 11713 8527 11747
rect 8585 11713 8619 11747
rect 8769 11713 8803 11747
rect 11529 11713 11563 11747
rect 11621 11713 11655 11747
rect 12081 11713 12115 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 12725 11713 12759 11747
rect 14841 11713 14875 11747
rect 17233 11713 17267 11747
rect 2697 11645 2731 11679
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 6101 11645 6135 11679
rect 8861 11645 8895 11679
rect 13001 11645 13035 11679
rect 13093 11645 13127 11679
rect 15025 11645 15059 11679
rect 4353 11577 4387 11611
rect 4445 11577 4479 11611
rect 5181 11577 5215 11611
rect 11897 11577 11931 11611
rect 17417 11577 17451 11611
rect 4077 11509 4111 11543
rect 7757 11509 7791 11543
rect 11989 11509 12023 11543
rect 12817 11509 12851 11543
rect 10793 11305 10827 11339
rect 12173 11305 12207 11339
rect 12817 11305 12851 11339
rect 17417 11305 17451 11339
rect 9045 11169 9079 11203
rect 15945 11169 15979 11203
rect 1409 11101 1443 11135
rect 12357 11101 12391 11135
rect 12449 11101 12483 11135
rect 12577 11101 12611 11135
rect 12909 11101 12943 11135
rect 15669 11101 15703 11135
rect 9321 11033 9355 11067
rect 12173 11033 12207 11067
rect 1593 10965 1627 10999
rect 2513 10761 2547 10795
rect 5181 10761 5215 10795
rect 5733 10761 5767 10795
rect 7113 10761 7147 10795
rect 10057 10761 10091 10795
rect 13185 10761 13219 10795
rect 14565 10761 14599 10795
rect 16129 10761 16163 10795
rect 17233 10761 17267 10795
rect 8769 10693 8803 10727
rect 10701 10693 10735 10727
rect 2605 10625 2639 10659
rect 4169 10625 4203 10659
rect 4261 10625 4295 10659
rect 4353 10625 4387 10659
rect 4537 10625 4571 10659
rect 4813 10625 4847 10659
rect 5395 10625 5429 10659
rect 5549 10625 5583 10659
rect 5825 10625 5859 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 7297 10625 7331 10659
rect 7757 10625 7791 10659
rect 7849 10625 7883 10659
rect 10793 10625 10827 10659
rect 11989 10625 12023 10659
rect 13001 10625 13035 10659
rect 13277 10625 13311 10659
rect 13369 10625 13403 10659
rect 13644 10625 13678 10659
rect 13737 10625 13771 10659
rect 14289 10625 14323 10659
rect 14933 10625 14967 10659
rect 17141 10625 17175 10659
rect 17417 10625 17451 10659
rect 2697 10557 2731 10591
rect 4629 10557 4663 10591
rect 4997 10557 5031 10591
rect 6561 10557 6595 10591
rect 6653 10557 6687 10591
rect 7481 10557 7515 10591
rect 13829 10557 13863 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 16221 10557 16255 10591
rect 16313 10557 16347 10591
rect 7389 10489 7423 10523
rect 13921 10489 13955 10523
rect 16957 10489 16991 10523
rect 2145 10421 2179 10455
rect 3893 10421 3927 10455
rect 12081 10421 12115 10455
rect 13001 10421 13035 10455
rect 15761 10421 15795 10455
rect 5273 10217 5307 10251
rect 8309 10217 8343 10251
rect 10977 10217 11011 10251
rect 17325 10217 17359 10251
rect 3801 10149 3835 10183
rect 1409 10081 1443 10115
rect 11437 10081 11471 10115
rect 11621 10081 11655 10115
rect 15853 10081 15887 10115
rect 3433 10013 3467 10047
rect 4077 10013 4111 10047
rect 4445 10013 4479 10047
rect 5198 10013 5232 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 6101 10013 6135 10047
rect 8125 10013 8159 10047
rect 8218 10013 8252 10047
rect 11805 10013 11839 10047
rect 15577 10013 15611 10047
rect 1685 9945 1719 9979
rect 3341 9945 3375 9979
rect 3801 9945 3835 9979
rect 4353 9945 4387 9979
rect 3157 9877 3191 9911
rect 3985 9877 4019 9911
rect 5733 9877 5767 9911
rect 11345 9877 11379 9911
rect 13093 9877 13127 9911
rect 6837 9673 6871 9707
rect 11069 9673 11103 9707
rect 8125 9605 8159 9639
rect 9505 9605 9539 9639
rect 9781 9605 9815 9639
rect 13461 9605 13495 9639
rect 16773 9605 16807 9639
rect 9137 9537 9171 9571
rect 9597 9537 9631 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 10885 9537 10919 9571
rect 11805 9537 11839 9571
rect 13553 9537 13587 9571
rect 14749 9537 14783 9571
rect 16865 9537 16899 9571
rect 17417 9537 17451 9571
rect 9045 9469 9079 9503
rect 9229 9469 9263 9503
rect 9321 9469 9355 9503
rect 10333 9469 10367 9503
rect 10793 9469 10827 9503
rect 11161 9469 11195 9503
rect 11253 9469 11287 9503
rect 12817 9469 12851 9503
rect 14841 9469 14875 9503
rect 15025 9469 15059 9503
rect 9597 9401 9631 9435
rect 13185 9401 13219 9435
rect 14381 9401 14415 9435
rect 17233 9401 17267 9435
rect 10057 9333 10091 9367
rect 13277 9333 13311 9367
rect 5825 9129 5859 9163
rect 13369 9129 13403 9163
rect 7297 9061 7331 9095
rect 12725 9061 12759 9095
rect 5733 8993 5767 9027
rect 5825 8993 5859 9027
rect 6929 8993 6963 9027
rect 7573 8993 7607 9027
rect 7665 8993 7699 9027
rect 7849 8993 7883 9027
rect 8033 8993 8067 9027
rect 12817 8993 12851 9027
rect 13185 8993 13219 9027
rect 15393 8993 15427 9027
rect 16589 8993 16623 9027
rect 3893 8925 3927 8959
rect 3986 8925 4020 8959
rect 5641 8925 5675 8959
rect 6837 8925 6871 8959
rect 7021 8925 7055 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 7941 8925 7975 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 8493 8925 8527 8959
rect 8677 8925 8711 8959
rect 12633 8925 12667 8959
rect 12909 8925 12943 8959
rect 13461 8925 13495 8959
rect 15117 8925 15151 8959
rect 16405 8925 16439 8959
rect 6009 8857 6043 8891
rect 7481 8857 7515 8891
rect 8585 8857 8619 8891
rect 13185 8857 13219 8891
rect 4261 8789 4295 8823
rect 13093 8789 13127 8823
rect 14749 8789 14783 8823
rect 15209 8789 15243 8823
rect 16037 8789 16071 8823
rect 16497 8789 16531 8823
rect 3341 8585 3375 8619
rect 6009 8585 6043 8619
rect 11897 8585 11931 8619
rect 13369 8585 13403 8619
rect 3617 8517 3651 8551
rect 13461 8517 13495 8551
rect 13645 8517 13679 8551
rect 3157 8449 3191 8483
rect 3433 8449 3467 8483
rect 3831 8449 3865 8483
rect 3985 8449 4019 8483
rect 4077 8449 4111 8483
rect 4261 8449 4295 8483
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 5272 8449 5306 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 7665 8449 7699 8483
rect 7941 8449 7975 8483
rect 8033 8449 8067 8483
rect 11529 8449 11563 8483
rect 11622 8449 11656 8483
rect 12817 8449 12851 8483
rect 13001 8449 13035 8483
rect 13093 8449 13127 8483
rect 13553 8449 13587 8483
rect 13920 8449 13954 8483
rect 14013 8449 14047 8483
rect 14472 8449 14506 8483
rect 14565 8449 14599 8483
rect 2881 8381 2915 8415
rect 5641 8381 5675 8415
rect 6377 8381 6411 8415
rect 6469 8381 6503 8415
rect 7757 8381 7791 8415
rect 13185 8381 13219 8415
rect 14197 8381 14231 8415
rect 6929 8313 6963 8347
rect 12633 8313 12667 8347
rect 13461 8313 13495 8347
rect 1409 8245 1443 8279
rect 7481 8245 7515 8279
rect 8217 8245 8251 8279
rect 1409 8041 1443 8075
rect 12265 8041 12299 8075
rect 17371 8041 17405 8075
rect 4261 7973 4295 8007
rect 10701 7973 10735 8007
rect 7113 7905 7147 7939
rect 10793 7905 10827 7939
rect 15945 7905 15979 7939
rect 1593 7837 1627 7871
rect 1869 7837 1903 7871
rect 3893 7837 3927 7871
rect 3986 7837 4020 7871
rect 6929 7837 6963 7871
rect 7481 7837 7515 7871
rect 8033 7837 8067 7871
rect 10333 7837 10367 7871
rect 12081 7837 12115 7871
rect 12174 7837 12208 7871
rect 15577 7837 15611 7871
rect 10517 7769 10551 7803
rect 1685 7701 1719 7735
rect 10057 7701 10091 7735
rect 10425 7701 10459 7735
rect 1409 7497 1443 7531
rect 8217 7497 8251 7531
rect 16037 7497 16071 7531
rect 16773 7497 16807 7531
rect 9597 7429 9631 7463
rect 11345 7429 11379 7463
rect 14565 7429 14599 7463
rect 16221 7429 16255 7463
rect 3157 7361 3191 7395
rect 8125 7361 8159 7395
rect 9045 7361 9079 7395
rect 9137 7361 9171 7395
rect 9321 7361 9355 7395
rect 14289 7361 14323 7395
rect 16313 7361 16347 7395
rect 16865 7361 16899 7395
rect 2881 7293 2915 7327
rect 8861 7157 8895 7191
rect 2605 6817 2639 6851
rect 4445 6817 4479 6851
rect 5733 6817 5767 6851
rect 8125 6817 8159 6851
rect 8585 6817 8619 6851
rect 9045 6817 9079 6851
rect 10701 6817 10735 6851
rect 12357 6817 12391 6851
rect 12817 6817 12851 6851
rect 2697 6749 2731 6783
rect 4353 6749 4387 6783
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 6653 6749 6687 6783
rect 8493 6749 8527 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 10793 6749 10827 6783
rect 12449 6749 12483 6783
rect 6101 6681 6135 6715
rect 6377 6681 6411 6715
rect 6469 6681 6503 6715
rect 3157 6409 3191 6443
rect 7481 6409 7515 6443
rect 7573 6409 7607 6443
rect 11345 6341 11379 6375
rect 11805 6341 11839 6375
rect 11989 6341 12023 6375
rect 13093 6341 13127 6375
rect 13553 6341 13587 6375
rect 4905 6273 4939 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 5917 6273 5951 6307
rect 6837 6273 6871 6307
rect 6929 6273 6963 6307
rect 7665 6273 7699 6307
rect 11069 6273 11103 6307
rect 11161 6273 11195 6307
rect 12633 6273 12667 6307
rect 12725 6273 12759 6307
rect 12817 6273 12851 6307
rect 4629 6205 4663 6239
rect 5181 6205 5215 6239
rect 7021 6205 7055 6239
rect 7113 6205 7147 6239
rect 7297 6205 7331 6239
rect 12357 6205 12391 6239
rect 13277 6205 13311 6239
rect 15301 6205 15335 6239
rect 5825 6137 5859 6171
rect 6653 6069 6687 6103
rect 7389 6069 7423 6103
rect 11345 6069 11379 6103
rect 11621 6069 11655 6103
rect 11805 6069 11839 6103
rect 12449 6069 12483 6103
rect 3985 5865 4019 5899
rect 14565 5865 14599 5899
rect 5733 5729 5767 5763
rect 9597 5729 9631 5763
rect 9873 5729 9907 5763
rect 4077 5661 4111 5695
rect 5917 5661 5951 5695
rect 9505 5661 9539 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 14657 5661 14691 5695
rect 6101 5525 6135 5559
rect 11713 5525 11747 5559
rect 6837 5321 6871 5355
rect 8401 5321 8435 5355
rect 10517 5321 10551 5355
rect 12541 5321 12575 5355
rect 12449 5253 12483 5287
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7021 5185 7055 5219
rect 8217 5185 8251 5219
rect 8309 5185 8343 5219
rect 8677 5185 8711 5219
rect 10333 5185 10367 5219
rect 10425 5185 10459 5219
rect 10793 5185 10827 5219
rect 12357 5185 12391 5219
rect 7113 5117 7147 5151
rect 12817 5117 12851 5151
rect 10701 5049 10735 5083
rect 12725 5049 12759 5083
rect 6377 4981 6411 5015
rect 7941 4981 7975 5015
rect 8585 4981 8619 5015
rect 10057 4981 10091 5015
rect 12081 4981 12115 5015
rect 12338 4777 12372 4811
rect 13829 4777 13863 4811
rect 5181 4641 5215 4675
rect 7205 4641 7239 4675
rect 9873 4641 9907 4675
rect 12081 4641 12115 4675
rect 8401 4573 8435 4607
rect 11897 4573 11931 4607
rect 14289 4573 14323 4607
rect 6929 4505 6963 4539
rect 10149 4505 10183 4539
rect 14197 4505 14231 4539
rect 8493 4437 8527 4471
rect 11069 4233 11103 4267
rect 7665 4165 7699 4199
rect 6469 4097 6503 4131
rect 6561 4097 6595 4131
rect 7389 4097 7423 4131
rect 9413 4097 9447 4131
rect 11161 4097 11195 4131
rect 16589 3553 16623 3587
rect 17417 3485 17451 3519
<< metal1 >>
rect 1104 18522 17756 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 17756 18522
rect 1104 18448 17756 18470
rect 7190 18368 7196 18420
rect 7248 18368 7254 18420
rect 7834 18368 7840 18420
rect 7892 18368 7898 18420
rect 8478 18368 8484 18420
rect 8536 18368 8542 18420
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 11698 18368 11704 18420
rect 11756 18368 11762 18420
rect 12986 18368 12992 18420
rect 13044 18368 13050 18420
rect 10502 18300 10508 18352
rect 10560 18300 10566 18352
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 3878 18272 3884 18284
rect 2363 18244 3884 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 6086 18232 6092 18284
rect 6144 18232 6150 18284
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7098 18272 7104 18284
rect 6871 18244 7104 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 7098 18232 7104 18244
rect 7156 18272 7162 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7156 18244 7389 18272
rect 7156 18232 7162 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7800 18244 8033 18272
rect 7800 18232 7806 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8021 18235 8079 18241
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 9306 18232 9312 18284
rect 9364 18232 9370 18284
rect 9950 18232 9956 18284
rect 10008 18232 10014 18284
rect 10870 18232 10876 18284
rect 10928 18272 10934 18284
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 10928 18244 11069 18272
rect 10928 18232 10934 18244
rect 11057 18241 11069 18244
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 11882 18232 11888 18284
rect 11940 18232 11946 18284
rect 12342 18232 12348 18284
rect 12400 18232 12406 18284
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 13188 18204 13216 18235
rect 13630 18232 13636 18284
rect 13688 18232 13694 18284
rect 13906 18204 13912 18216
rect 13188 18176 13912 18204
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 10686 18096 10692 18148
rect 10744 18096 10750 18148
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2409 18071 2467 18077
rect 2409 18068 2421 18071
rect 2188 18040 2421 18068
rect 2188 18028 2194 18040
rect 2409 18037 2421 18040
rect 2455 18037 2467 18071
rect 2409 18031 2467 18037
rect 4522 18028 4528 18080
rect 4580 18068 4586 18080
rect 5905 18071 5963 18077
rect 5905 18068 5917 18071
rect 4580 18040 5917 18068
rect 4580 18028 4586 18040
rect 5905 18037 5917 18040
rect 5951 18037 5963 18071
rect 5905 18031 5963 18037
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6052 18040 6377 18068
rect 6052 18028 6058 18040
rect 6365 18037 6377 18040
rect 6411 18037 6423 18071
rect 6365 18031 6423 18037
rect 6733 18071 6791 18077
rect 6733 18037 6745 18071
rect 6779 18068 6791 18071
rect 6914 18068 6920 18080
rect 6779 18040 6920 18068
rect 6779 18037 6791 18040
rect 6733 18031 6791 18037
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 9769 18071 9827 18077
rect 9769 18068 9781 18071
rect 9732 18040 9781 18068
rect 9732 18028 9738 18040
rect 9769 18037 9781 18040
rect 9815 18037 9827 18071
rect 9769 18031 9827 18037
rect 11241 18071 11299 18077
rect 11241 18037 11253 18071
rect 11287 18068 11299 18071
rect 11514 18068 11520 18080
rect 11287 18040 11520 18068
rect 11287 18037 11299 18040
rect 11241 18031 11299 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 12526 18028 12532 18080
rect 12584 18028 12590 18080
rect 13814 18028 13820 18080
rect 13872 18028 13878 18080
rect 1104 17978 17756 18000
rect 1104 17926 2350 17978
rect 2402 17926 2414 17978
rect 2466 17926 2478 17978
rect 2530 17926 2542 17978
rect 2594 17926 2606 17978
rect 2658 17926 17756 17978
rect 1104 17904 17756 17926
rect 7098 17824 7104 17876
rect 7156 17824 7162 17876
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 11940 17836 12081 17864
rect 11940 17824 11946 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 13906 17824 13912 17876
rect 13964 17824 13970 17876
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 2774 17728 2780 17740
rect 1443 17700 2780 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 2774 17688 2780 17700
rect 2832 17728 2838 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 2832 17700 3801 17728
rect 2832 17688 2838 17700
rect 3789 17697 3801 17700
rect 3835 17728 3847 17731
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 3835 17700 5764 17728
rect 3835 17697 3847 17700
rect 3789 17691 3847 17697
rect 1762 17620 1768 17672
rect 1820 17620 1826 17672
rect 4154 17620 4160 17672
rect 4212 17620 4218 17672
rect 5736 17669 5764 17700
rect 12176 17700 14657 17728
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17660 5779 17663
rect 6362 17660 6368 17672
rect 5767 17632 6368 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 6362 17620 6368 17632
rect 6420 17660 6426 17672
rect 12176 17669 12204 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 6420 17632 7389 17660
rect 6420 17620 6426 17632
rect 7377 17629 7389 17632
rect 7423 17629 7435 17663
rect 7377 17623 7435 17629
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17660 9275 17663
rect 10689 17663 10747 17669
rect 10689 17660 10701 17663
rect 9263 17632 10701 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 10689 17629 10701 17632
rect 10735 17660 10747 17663
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 10735 17632 12173 17660
rect 10735 17629 10747 17632
rect 10689 17623 10747 17629
rect 11072 17604 11100 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 14274 17620 14280 17672
rect 14332 17620 14338 17672
rect 14660 17660 14688 17691
rect 15654 17660 15660 17672
rect 14660 17632 15660 17660
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 2130 17552 2136 17604
rect 2188 17552 2194 17604
rect 5994 17601 6000 17604
rect 5988 17592 6000 17601
rect 4448 17564 4554 17592
rect 5955 17564 6000 17592
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 3191 17527 3249 17533
rect 3191 17524 3203 17527
rect 2556 17496 3203 17524
rect 2556 17484 2562 17496
rect 3191 17493 3203 17496
rect 3237 17493 3249 17527
rect 3191 17487 3249 17493
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4448 17524 4476 17564
rect 5988 17555 6000 17564
rect 5994 17552 6000 17555
rect 6052 17552 6058 17604
rect 7644 17595 7702 17601
rect 7644 17561 7656 17595
rect 7690 17592 7702 17595
rect 7834 17592 7840 17604
rect 7690 17564 7840 17592
rect 7690 17561 7702 17564
rect 7644 17555 7702 17561
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 9490 17601 9496 17604
rect 9484 17555 9496 17601
rect 9490 17552 9496 17555
rect 9548 17552 9554 17604
rect 10962 17601 10968 17604
rect 10956 17555 10968 17601
rect 10962 17552 10968 17555
rect 11020 17552 11026 17604
rect 11054 17552 11060 17604
rect 11112 17552 11118 17604
rect 14918 17601 14924 17604
rect 12437 17595 12495 17601
rect 12437 17561 12449 17595
rect 12483 17561 12495 17595
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 13662 17564 14197 17592
rect 12437 17555 12495 17561
rect 14185 17561 14197 17564
rect 14231 17561 14243 17595
rect 14185 17555 14243 17561
rect 14912 17555 14924 17601
rect 4120 17496 4476 17524
rect 4120 17484 4126 17496
rect 4614 17484 4620 17536
rect 4672 17524 4678 17536
rect 5583 17527 5641 17533
rect 5583 17524 5595 17527
rect 4672 17496 5595 17524
rect 4672 17484 4678 17496
rect 5583 17493 5595 17496
rect 5629 17524 5641 17527
rect 6454 17524 6460 17536
rect 5629 17496 6460 17524
rect 5629 17493 5641 17496
rect 5583 17487 5641 17493
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8662 17524 8668 17536
rect 8352 17496 8668 17524
rect 8352 17484 8358 17496
rect 8662 17484 8668 17496
rect 8720 17524 8726 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8720 17496 8769 17524
rect 8720 17484 8726 17496
rect 8757 17493 8769 17496
rect 8803 17493 8815 17527
rect 8757 17487 8815 17493
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 12452 17524 12480 17555
rect 14918 17552 14924 17555
rect 14976 17552 14982 17604
rect 10652 17496 12480 17524
rect 10652 17484 10658 17496
rect 16022 17484 16028 17536
rect 16080 17484 16086 17536
rect 1104 17434 17756 17456
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 17756 17434
rect 1104 17360 17756 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 2041 17323 2099 17329
rect 2041 17320 2053 17323
rect 1820 17292 2053 17320
rect 1820 17280 1826 17292
rect 2041 17289 2053 17292
rect 2087 17289 2099 17323
rect 2041 17283 2099 17289
rect 2498 17280 2504 17332
rect 2556 17280 2562 17332
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4062 17320 4068 17332
rect 4019 17292 4068 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4154 17280 4160 17332
rect 4212 17280 4218 17332
rect 4522 17280 4528 17332
rect 4580 17280 4586 17332
rect 4614 17280 4620 17332
rect 4672 17280 4678 17332
rect 7742 17280 7748 17332
rect 7800 17280 7806 17332
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 11020 17292 11529 17320
rect 11020 17280 11026 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17320 13783 17323
rect 13906 17320 13912 17332
rect 13771 17292 13912 17320
rect 13771 17289 13783 17292
rect 13725 17283 13783 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 2516 17252 2544 17280
rect 5902 17252 5908 17264
rect 2516 17224 5908 17252
rect 5902 17212 5908 17224
rect 5960 17212 5966 17264
rect 9416 17224 9812 17252
rect 9416 17196 9444 17224
rect 2222 17144 2228 17196
rect 2280 17184 2286 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2280 17156 2421 17184
rect 2280 17144 2286 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 3878 17144 3884 17196
rect 3936 17144 3942 17196
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6638 17193 6644 17196
rect 6632 17147 6644 17193
rect 6638 17144 6644 17147
rect 6696 17144 6702 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 6972 17156 7972 17184
rect 6972 17144 6978 17156
rect 2130 17076 2136 17128
rect 2188 17116 2194 17128
rect 2685 17119 2743 17125
rect 2685 17116 2697 17119
rect 2188 17088 2697 17116
rect 2188 17076 2194 17088
rect 2685 17085 2697 17088
rect 2731 17116 2743 17119
rect 4706 17116 4712 17128
rect 2731 17088 4712 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7944 17116 7972 17156
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 8294 17144 8300 17196
rect 8352 17144 8358 17196
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17184 9367 17187
rect 9398 17184 9404 17196
rect 9355 17156 9404 17184
rect 9355 17153 9367 17156
rect 9309 17147 9367 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9582 17184 9588 17196
rect 9508 17156 9588 17184
rect 8202 17116 8208 17128
rect 7944 17088 8208 17116
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 9508 17125 9536 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 9784 17193 9812 17224
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 9950 17144 9956 17196
rect 10008 17144 10014 17196
rect 10594 17144 10600 17196
rect 10652 17144 10658 17196
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11940 17156 11989 17184
rect 11940 17144 11946 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 13817 17187 13875 17193
rect 13817 17153 13829 17187
rect 13863 17184 13875 17187
rect 13998 17184 14004 17196
rect 13863 17156 14004 17184
rect 13863 17153 13875 17156
rect 13817 17147 13875 17153
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 9493 17079 9551 17085
rect 9600 17088 10517 17116
rect 9401 17051 9459 17057
rect 9401 17017 9413 17051
rect 9447 17048 9459 17051
rect 9600 17048 9628 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 13372 17116 13400 17147
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 14332 17156 16313 17184
rect 14332 17144 14338 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 13633 17119 13691 17125
rect 13633 17116 13645 17119
rect 13372 17088 13645 17116
rect 10505 17079 10563 17085
rect 13633 17085 13645 17088
rect 13679 17085 13691 17119
rect 13633 17079 13691 17085
rect 9447 17020 9628 17048
rect 9677 17051 9735 17057
rect 9447 17017 9459 17020
rect 9401 17011 9459 17017
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 9723 17020 9873 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 13648 17048 13676 17079
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 17000 17088 17141 17116
rect 17000 17076 17006 17088
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 13814 17048 13820 17060
rect 9861 17011 9919 17017
rect 12406 17020 13584 17048
rect 13648 17020 13820 17048
rect 9490 16940 9496 16992
rect 9548 16940 9554 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12406 16980 12434 17020
rect 11940 16952 12434 16980
rect 11940 16940 11946 16952
rect 13078 16940 13084 16992
rect 13136 16980 13142 16992
rect 13265 16983 13323 16989
rect 13265 16980 13277 16983
rect 13136 16952 13277 16980
rect 13136 16940 13142 16952
rect 13265 16949 13277 16952
rect 13311 16949 13323 16983
rect 13556 16980 13584 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 15102 17048 15108 17060
rect 14016 17020 15108 17048
rect 14016 16980 14044 17020
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 16758 17008 16764 17060
rect 16816 17048 16822 17060
rect 17236 17048 17264 17079
rect 16816 17020 17264 17048
rect 16816 17008 16822 17020
rect 13556 16952 14044 16980
rect 13265 16943 13323 16949
rect 14090 16940 14096 16992
rect 14148 16980 14154 16992
rect 14185 16983 14243 16989
rect 14185 16980 14197 16983
rect 14148 16952 14197 16980
rect 14148 16940 14154 16952
rect 14185 16949 14197 16952
rect 14231 16949 14243 16983
rect 14185 16943 14243 16949
rect 16393 16983 16451 16989
rect 16393 16949 16405 16983
rect 16439 16980 16451 16983
rect 16574 16980 16580 16992
rect 16439 16952 16580 16980
rect 16439 16949 16451 16952
rect 16393 16943 16451 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 1104 16890 17756 16912
rect 1104 16838 2350 16890
rect 2402 16838 2414 16890
rect 2466 16838 2478 16890
rect 2530 16838 2542 16890
rect 2594 16838 2606 16890
rect 2658 16838 17756 16890
rect 1104 16816 17756 16838
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 6638 16776 6644 16788
rect 6595 16748 6644 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 6914 16736 6920 16788
rect 6972 16736 6978 16788
rect 8202 16736 8208 16788
rect 8260 16776 8266 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 8260 16748 9413 16776
rect 8260 16736 8266 16748
rect 9401 16745 9413 16748
rect 9447 16776 9459 16779
rect 11882 16776 11888 16788
rect 9447 16748 11888 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 10962 16708 10968 16720
rect 4764 16680 10968 16708
rect 4764 16668 4770 16680
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16640 7067 16643
rect 7742 16640 7748 16652
rect 7055 16612 7748 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 9490 16600 9496 16652
rect 9548 16640 9554 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9548 16612 9781 16640
rect 9548 16600 9554 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 15654 16600 15660 16652
rect 15712 16600 15718 16652
rect 15933 16643 15991 16649
rect 15933 16609 15945 16643
rect 15979 16640 15991 16643
rect 16666 16640 16672 16652
rect 15979 16612 16672 16640
rect 15979 16609 15991 16612
rect 15933 16603 15991 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 6730 16532 6736 16584
rect 6788 16532 6794 16584
rect 9585 16575 9643 16581
rect 9585 16541 9597 16575
rect 9631 16572 9643 16575
rect 9674 16572 9680 16584
rect 9631 16544 9680 16572
rect 9631 16541 9643 16544
rect 9585 16535 9643 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 16574 16464 16580 16516
rect 16632 16464 16638 16516
rect 14182 16396 14188 16448
rect 14240 16436 14246 16448
rect 16942 16436 16948 16448
rect 14240 16408 16948 16436
rect 14240 16396 14246 16408
rect 16942 16396 16948 16408
rect 17000 16436 17006 16448
rect 17405 16439 17463 16445
rect 17405 16436 17417 16439
rect 17000 16408 17417 16436
rect 17000 16396 17006 16408
rect 17405 16405 17417 16408
rect 17451 16405 17463 16439
rect 17405 16399 17463 16405
rect 1104 16346 17756 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 17756 16346
rect 1104 16272 17756 16294
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14829 16235 14887 16241
rect 14829 16232 14841 16235
rect 14047 16204 14841 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14829 16201 14841 16204
rect 14875 16201 14887 16235
rect 14829 16195 14887 16201
rect 14918 16192 14924 16244
rect 14976 16192 14982 16244
rect 14090 16124 14096 16176
rect 14148 16124 14154 16176
rect 2777 16099 2835 16105
rect 2777 16065 2789 16099
rect 2823 16096 2835 16099
rect 3878 16096 3884 16108
rect 2823 16068 3884 16096
rect 2823 16065 2835 16068
rect 2777 16059 2835 16065
rect 3878 16056 3884 16068
rect 3936 16096 3942 16108
rect 5442 16096 5448 16108
rect 3936 16068 5448 16096
rect 3936 16056 3942 16068
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 13832 15960 13860 16059
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14550 16096 14556 16108
rect 14323 16068 14556 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 15102 16056 15108 16108
rect 15160 16056 15166 16108
rect 15289 16099 15347 16105
rect 15289 16065 15301 16099
rect 15335 16096 15347 16099
rect 16022 16096 16028 16108
rect 15335 16068 16028 16096
rect 15335 16065 15347 16068
rect 15289 16059 15347 16065
rect 16022 16056 16028 16068
rect 16080 16096 16086 16108
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 16080 16068 17233 16096
rect 16080 16056 16086 16068
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 14090 15988 14096 16040
rect 14148 16028 14154 16040
rect 14200 16028 14228 16056
rect 14148 16000 14228 16028
rect 14148 15988 14154 16000
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 14458 15960 14464 15972
rect 13832 15932 14464 15960
rect 14458 15920 14464 15932
rect 14516 15920 14522 15972
rect 2682 15852 2688 15904
rect 2740 15852 2746 15904
rect 11330 15852 11336 15904
rect 11388 15892 11394 15904
rect 12250 15892 12256 15904
rect 11388 15864 12256 15892
rect 11388 15852 11394 15864
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 1104 15802 17756 15824
rect 1104 15750 2350 15802
rect 2402 15750 2414 15802
rect 2466 15750 2478 15802
rect 2530 15750 2542 15802
rect 2594 15750 2606 15802
rect 2658 15750 17756 15802
rect 1104 15728 17756 15750
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3375 15691 3433 15697
rect 3375 15688 3387 15691
rect 2924 15660 3387 15688
rect 2924 15648 2930 15660
rect 3375 15657 3387 15660
rect 3421 15688 3433 15691
rect 3421 15660 5580 15688
rect 3421 15657 3433 15660
rect 3375 15651 3433 15657
rect 5552 15620 5580 15660
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6788 15660 6929 15688
rect 6788 15648 6794 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 8018 15688 8024 15700
rect 7699 15660 8024 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 11974 15688 11980 15700
rect 10100 15660 11980 15688
rect 10100 15648 10106 15660
rect 11974 15648 11980 15660
rect 12032 15688 12038 15700
rect 12032 15660 12434 15688
rect 12032 15648 12038 15660
rect 7926 15620 7932 15632
rect 5552 15592 7932 15620
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 12406 15620 12434 15660
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 13630 15688 13636 15700
rect 12584 15660 13636 15688
rect 12584 15648 12590 15660
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 13906 15688 13912 15700
rect 13863 15660 13912 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 13998 15620 14004 15632
rect 12406 15592 14004 15620
rect 13998 15580 14004 15592
rect 14056 15580 14062 15632
rect 2774 15552 2780 15564
rect 1596 15524 2780 15552
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 1596 15493 1624 15524
rect 2774 15512 2780 15524
rect 2832 15552 2838 15564
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 2832 15524 3801 15552
rect 2832 15512 2838 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 5902 15512 5908 15564
rect 5960 15552 5966 15564
rect 5960 15524 7144 15552
rect 5960 15512 5966 15524
rect 1581 15487 1639 15493
rect 1581 15484 1593 15487
rect 1452 15456 1593 15484
rect 1452 15444 1458 15456
rect 1581 15453 1593 15456
rect 1627 15453 1639 15487
rect 1581 15447 1639 15453
rect 1946 15444 1952 15496
rect 2004 15444 2010 15496
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5500 15456 5825 15484
rect 5500 15444 5506 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 5813 15447 5871 15453
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 6454 15493 6460 15496
rect 6421 15487 6460 15493
rect 6421 15453 6433 15487
rect 6421 15447 6460 15453
rect 6454 15444 6460 15447
rect 6512 15444 6518 15496
rect 6730 15444 6736 15496
rect 6788 15493 6794 15496
rect 6788 15487 6815 15493
rect 6803 15453 6815 15487
rect 6788 15447 6815 15453
rect 6788 15444 6794 15447
rect 6914 15444 6920 15496
rect 6972 15444 6978 15496
rect 7006 15444 7012 15496
rect 7064 15444 7070 15496
rect 7116 15493 7144 15524
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 8205 15555 8263 15561
rect 8205 15552 8217 15555
rect 7340 15524 8217 15552
rect 7340 15512 7346 15524
rect 8205 15521 8217 15524
rect 8251 15521 8263 15555
rect 8205 15515 8263 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 7558 15493 7564 15496
rect 7102 15487 7160 15493
rect 7102 15453 7114 15487
rect 7148 15453 7160 15487
rect 7102 15447 7160 15453
rect 7515 15487 7564 15493
rect 7515 15453 7527 15487
rect 7561 15453 7564 15487
rect 7515 15447 7564 15453
rect 7558 15444 7564 15447
rect 7616 15444 7622 15496
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 8110 15484 8116 15496
rect 7708 15456 8116 15484
rect 7708 15444 7714 15456
rect 8110 15444 8116 15456
rect 8168 15484 8174 15496
rect 8312 15484 8340 15515
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 12158 15512 12164 15564
rect 12216 15512 12222 15564
rect 12529 15555 12587 15561
rect 12529 15552 12541 15555
rect 12406 15524 12541 15552
rect 8168 15456 8340 15484
rect 8168 15444 8174 15456
rect 11330 15444 11336 15496
rect 11388 15444 11394 15496
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 11900 15484 12020 15486
rect 12406 15484 12434 15524
rect 12529 15521 12541 15524
rect 12575 15552 12587 15555
rect 12575 15524 13584 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13556 15496 13584 15524
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 15933 15555 15991 15561
rect 15933 15552 15945 15555
rect 15712 15524 15945 15552
rect 15712 15512 15718 15524
rect 15933 15521 15945 15524
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 11572 15458 12434 15484
rect 11572 15456 11928 15458
rect 11992 15456 12434 15458
rect 12544 15456 13001 15484
rect 11572 15444 11578 15456
rect 2682 15376 2688 15428
rect 2740 15376 2746 15428
rect 4065 15419 4123 15425
rect 4065 15385 4077 15419
rect 4111 15416 4123 15419
rect 4338 15416 4344 15428
rect 4111 15388 4344 15416
rect 4111 15385 4123 15388
rect 4065 15379 4123 15385
rect 4338 15376 4344 15388
rect 4396 15376 4402 15428
rect 5721 15419 5779 15425
rect 5721 15416 5733 15419
rect 5290 15388 5733 15416
rect 5721 15385 5733 15388
rect 5767 15385 5779 15419
rect 5721 15379 5779 15385
rect 6178 15376 6184 15428
rect 6236 15416 6242 15428
rect 6549 15419 6607 15425
rect 6549 15416 6561 15419
rect 6236 15388 6561 15416
rect 6236 15376 6242 15388
rect 6549 15385 6561 15388
rect 6595 15385 6607 15419
rect 6549 15379 6607 15385
rect 6641 15419 6699 15425
rect 6641 15385 6653 15419
rect 6687 15416 6699 15419
rect 6932 15416 6960 15444
rect 6687 15388 6960 15416
rect 7285 15419 7343 15425
rect 6687 15385 6699 15388
rect 6641 15379 6699 15385
rect 7285 15385 7297 15419
rect 7331 15385 7343 15419
rect 7285 15379 7343 15385
rect 7377 15419 7435 15425
rect 7377 15385 7389 15419
rect 7423 15416 7435 15419
rect 7423 15388 7788 15416
rect 7423 15385 7435 15388
rect 7377 15379 7435 15385
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 6822 15348 6828 15360
rect 5592 15320 6828 15348
rect 5592 15308 5598 15320
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7300 15348 7328 15379
rect 7466 15348 7472 15360
rect 7300 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 7760 15357 7788 15388
rect 9030 15376 9036 15428
rect 9088 15376 9094 15428
rect 9490 15376 9496 15428
rect 9548 15416 9554 15428
rect 10781 15419 10839 15425
rect 9548 15388 9614 15416
rect 9548 15376 9554 15388
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 10827 15388 11652 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 7745 15351 7803 15357
rect 7745 15317 7757 15351
rect 7791 15317 7803 15351
rect 7745 15311 7803 15317
rect 8018 15308 8024 15360
rect 8076 15348 8082 15360
rect 8113 15351 8171 15357
rect 8113 15348 8125 15351
rect 8076 15320 8125 15348
rect 8076 15308 8082 15320
rect 8113 15317 8125 15320
rect 8159 15317 8171 15351
rect 9048 15348 9076 15376
rect 9950 15348 9956 15360
rect 9048 15320 9956 15348
rect 8113 15311 8171 15317
rect 9950 15308 9956 15320
rect 10008 15308 10014 15360
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 11624 15357 11652 15388
rect 11974 15376 11980 15428
rect 12032 15376 12038 15428
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12544 15416 12572 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 12308 15388 12572 15416
rect 12308 15376 12314 15388
rect 12618 15376 12624 15428
rect 12676 15376 12682 15428
rect 13004 15416 13032 15447
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 13170 15444 13176 15496
rect 13228 15444 13234 15496
rect 13538 15444 13544 15496
rect 13596 15444 13602 15496
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13688 15456 14105 15484
rect 13688 15444 13694 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 17218 15484 17224 15496
rect 14323 15456 17224 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 13004 15388 13461 15416
rect 13449 15385 13461 15388
rect 13495 15416 13507 15419
rect 13722 15416 13728 15428
rect 13495 15388 13728 15416
rect 13495 15385 13507 15388
rect 13449 15379 13507 15385
rect 13722 15376 13728 15388
rect 13780 15376 13786 15428
rect 13817 15419 13875 15425
rect 13817 15385 13829 15419
rect 13863 15416 13875 15419
rect 14292 15416 14320 15447
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 13863 15388 14320 15416
rect 13863 15385 13875 15388
rect 13817 15379 13875 15385
rect 15838 15376 15844 15428
rect 15896 15416 15902 15428
rect 16178 15419 16236 15425
rect 16178 15416 16190 15419
rect 15896 15388 16190 15416
rect 15896 15376 15902 15388
rect 16178 15385 16190 15388
rect 16224 15385 16236 15419
rect 16178 15379 16236 15385
rect 11609 15351 11667 15357
rect 11609 15317 11621 15351
rect 11655 15317 11667 15351
rect 11609 15311 11667 15317
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12894 15348 12900 15360
rect 12115 15320 12900 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13262 15308 13268 15360
rect 13320 15348 13326 15360
rect 14185 15351 14243 15357
rect 14185 15348 14197 15351
rect 13320 15320 14197 15348
rect 13320 15308 13326 15320
rect 14185 15317 14197 15320
rect 14231 15317 14243 15351
rect 14185 15311 14243 15317
rect 17310 15308 17316 15360
rect 17368 15308 17374 15360
rect 1104 15258 17756 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 17756 15258
rect 1104 15184 17756 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 2225 15147 2283 15153
rect 2225 15144 2237 15147
rect 2004 15116 2237 15144
rect 2004 15104 2010 15116
rect 2225 15113 2237 15116
rect 2271 15113 2283 15147
rect 2225 15107 2283 15113
rect 2685 15147 2743 15153
rect 2685 15113 2697 15147
rect 2731 15144 2743 15147
rect 2866 15144 2872 15156
rect 2731 15116 2872 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4338 15104 4344 15156
rect 4396 15144 4402 15156
rect 4525 15147 4583 15153
rect 4525 15144 4537 15147
rect 4396 15116 4537 15144
rect 4396 15104 4402 15116
rect 4525 15113 4537 15116
rect 4571 15113 4583 15147
rect 4525 15107 4583 15113
rect 4985 15147 5043 15153
rect 4985 15113 4997 15147
rect 5031 15144 5043 15147
rect 5534 15144 5540 15156
rect 5031 15116 5540 15144
rect 5031 15113 5043 15116
rect 4985 15107 5043 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 6914 15104 6920 15156
rect 6972 15104 6978 15156
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 9398 15144 9404 15156
rect 7064 15116 9404 15144
rect 7064 15104 7070 15116
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 9490 15104 9496 15156
rect 9548 15104 9554 15156
rect 11330 15144 11336 15156
rect 10060 15116 11336 15144
rect 6730 15036 6736 15088
rect 6788 15076 6794 15088
rect 7558 15076 7564 15088
rect 6788 15048 7564 15076
rect 6788 15036 6794 15048
rect 7558 15036 7564 15048
rect 7616 15076 7622 15088
rect 7616 15048 7880 15076
rect 7616 15036 7622 15048
rect 842 14968 848 15020
rect 900 15008 906 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 900 14980 1409 15008
rect 900 14968 906 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 2222 14968 2228 15020
rect 2280 15008 2286 15020
rect 2593 15011 2651 15017
rect 2593 15008 2605 15011
rect 2280 14980 2605 15008
rect 2280 14968 2286 14980
rect 2593 14977 2605 14980
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4580 14980 4905 15008
rect 4580 14968 4586 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 6914 14968 6920 15020
rect 6972 15008 6978 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6972 14980 7297 15008
rect 6972 14968 6978 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7285 14971 7343 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7742 15008 7748 15020
rect 7423 14980 7748 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 2240 14872 2268 14968
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2372 14912 2881 14940
rect 2372 14900 2378 14912
rect 2869 14909 2881 14912
rect 2915 14940 2927 14943
rect 5169 14943 5227 14949
rect 2915 14912 4476 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 4448 14884 4476 14912
rect 5169 14909 5181 14943
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 1627 14844 2268 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 4430 14832 4436 14884
rect 4488 14872 4494 14884
rect 5184 14872 5212 14903
rect 5994 14900 6000 14952
rect 6052 14940 6058 14952
rect 6270 14940 6276 14952
rect 6052 14912 6276 14940
rect 6052 14900 6058 14912
rect 6270 14900 6276 14912
rect 6328 14940 6334 14952
rect 7006 14940 7012 14952
rect 6328 14912 7012 14940
rect 6328 14900 6334 14912
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7156 14912 7481 14940
rect 7156 14900 7162 14912
rect 7469 14909 7481 14912
rect 7515 14940 7527 14943
rect 7650 14940 7656 14952
rect 7515 14912 7656 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7852 14940 7880 15048
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 10060 15076 10088 15116
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11422 15104 11428 15156
rect 11480 15144 11486 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11480 15116 11897 15144
rect 11480 15104 11486 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 12158 15104 12164 15156
rect 12216 15104 12222 15156
rect 13078 15144 13084 15156
rect 12406 15116 13084 15144
rect 11609 15079 11667 15085
rect 11609 15076 11621 15079
rect 8168 15048 10088 15076
rect 8168 15036 8174 15048
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 9950 15008 9956 15020
rect 9631 14980 9956 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10060 15017 10088 15048
rect 10704 15048 11621 15076
rect 10704 15020 10732 15048
rect 11609 15045 11621 15048
rect 11655 15045 11667 15079
rect 11609 15039 11667 15045
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 12406 15076 12434 15116
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 14553 15147 14611 15153
rect 14553 15113 14565 15147
rect 14599 15144 14611 15147
rect 14734 15144 14740 15156
rect 14599 15116 14740 15144
rect 14599 15113 14611 15116
rect 14553 15107 14611 15113
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 15838 15104 15844 15156
rect 15896 15104 15902 15156
rect 12989 15079 13047 15085
rect 12989 15076 13001 15079
rect 12023 15048 12434 15076
rect 12544 15048 13001 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 10796 14980 11161 15008
rect 10796 14940 10824 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 14977 11851 15011
rect 12544 15008 12572 15048
rect 12989 15045 13001 15048
rect 13035 15076 13047 15079
rect 13262 15076 13268 15088
rect 13035 15048 13268 15076
rect 13035 15045 13047 15048
rect 12989 15039 13047 15045
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 11793 14971 11851 14977
rect 12084 14980 12572 15008
rect 12897 15011 12955 15017
rect 7852 14912 10824 14940
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 10980 14872 11008 14903
rect 11164 14884 11192 14971
rect 11808 14940 11836 14971
rect 12084 14940 12112 14980
rect 12897 14977 12909 15011
rect 12943 15008 12955 15011
rect 13078 15008 13084 15020
rect 12943 14980 13084 15008
rect 12943 14977 12955 14980
rect 12897 14971 12955 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 14366 14968 14372 15020
rect 14424 14968 14430 15020
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 11808 14912 12112 14940
rect 12176 14912 12449 14940
rect 4488 14844 11008 14872
rect 4488 14832 4494 14844
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 9950 14804 9956 14816
rect 5500 14776 9956 14804
rect 5500 14764 5506 14776
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10980 14804 11008 14844
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 12176 14872 12204 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13538 14940 13544 14952
rect 13219 14912 13544 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 11204 14844 12204 14872
rect 12452 14872 12480 14903
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 14568 14872 14596 14971
rect 16022 14968 16028 15020
rect 16080 14968 16086 15020
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 16114 14940 16120 14952
rect 15252 14912 16120 14940
rect 15252 14900 15258 14912
rect 16114 14900 16120 14912
rect 16172 14940 16178 14952
rect 16209 14943 16267 14949
rect 16209 14940 16221 14943
rect 16172 14912 16221 14940
rect 16172 14900 16178 14912
rect 16209 14909 16221 14912
rect 16255 14909 16267 14943
rect 16209 14903 16267 14909
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 17310 14940 17316 14952
rect 16347 14912 17316 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 14918 14872 14924 14884
rect 12452 14844 14924 14872
rect 11204 14832 11210 14844
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 12802 14804 12808 14816
rect 10980 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 1104 14714 17756 14736
rect 1104 14662 2350 14714
rect 2402 14662 2414 14714
rect 2466 14662 2478 14714
rect 2530 14662 2542 14714
rect 2594 14662 2606 14714
rect 2658 14662 17756 14714
rect 1104 14640 17756 14662
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6604 14572 6653 14600
rect 6604 14560 6610 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 6641 14563 6699 14569
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 17034 14600 17040 14612
rect 12952 14572 17040 14600
rect 12952 14560 12958 14572
rect 17034 14560 17040 14572
rect 17092 14600 17098 14612
rect 17221 14603 17279 14609
rect 17221 14600 17233 14603
rect 17092 14572 17233 14600
rect 17092 14560 17098 14572
rect 17221 14569 17233 14572
rect 17267 14569 17279 14603
rect 17221 14563 17279 14569
rect 6454 14492 6460 14544
rect 6512 14532 6518 14544
rect 7558 14532 7564 14544
rect 6512 14504 7564 14532
rect 6512 14492 6518 14504
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 7466 14464 7472 14476
rect 6236 14436 7472 14464
rect 6236 14424 6242 14436
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14396 2375 14399
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 2363 14368 4261 14396
rect 2363 14365 2375 14368
rect 2317 14359 2375 14365
rect 4249 14365 4261 14368
rect 4295 14396 4307 14399
rect 5442 14396 5448 14408
rect 4295 14368 5448 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 5994 14356 6000 14408
rect 6052 14356 6058 14408
rect 6086 14356 6092 14408
rect 6144 14396 6150 14408
rect 6288 14405 6316 14436
rect 7466 14424 7472 14436
rect 7524 14464 7530 14476
rect 12618 14464 12624 14476
rect 7524 14436 12624 14464
rect 7524 14424 7530 14436
rect 11348 14408 11376 14436
rect 12618 14424 12624 14436
rect 12676 14464 12682 14476
rect 14550 14464 14556 14476
rect 12676 14436 14556 14464
rect 12676 14424 12682 14436
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 6273 14399 6331 14405
rect 6144 14368 6189 14396
rect 6144 14356 6150 14368
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6503 14399 6561 14405
rect 6503 14365 6515 14399
rect 6549 14396 6561 14399
rect 6730 14396 6736 14408
rect 6549 14368 6736 14396
rect 6549 14365 6561 14368
rect 6503 14359 6561 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 17402 14356 17408 14408
rect 17460 14356 17466 14408
rect 6362 14288 6368 14340
rect 6420 14288 6426 14340
rect 2406 14220 2412 14272
rect 2464 14220 2470 14272
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 4304 14232 4353 14260
rect 4304 14220 4310 14232
rect 4341 14229 4353 14232
rect 4387 14229 4399 14263
rect 4341 14223 4399 14229
rect 1104 14170 17756 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 17756 14170
rect 1104 14096 17756 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1452 14028 3372 14056
rect 1452 14016 1458 14028
rect 2406 13948 2412 14000
rect 2464 13948 2470 14000
rect 3344 13932 3372 14028
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8444 14028 9045 14056
rect 8444 14016 8450 14028
rect 9033 14025 9045 14028
rect 9079 14056 9091 14059
rect 9306 14056 9312 14068
rect 9079 14028 9312 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 11241 14059 11299 14065
rect 11241 14025 11253 14059
rect 11287 14056 11299 14059
rect 11698 14056 11704 14068
rect 11287 14028 11704 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12529 14059 12587 14065
rect 12529 14025 12541 14059
rect 12575 14056 12587 14059
rect 12894 14056 12900 14068
rect 12575 14028 12900 14056
rect 12575 14025 12587 14028
rect 12529 14019 12587 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 14366 14016 14372 14068
rect 14424 14016 14430 14068
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 4246 13948 4252 14000
rect 4304 13948 4310 14000
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 10873 13991 10931 13997
rect 9456 13960 10640 13988
rect 9456 13948 9462 13960
rect 3326 13880 3332 13932
rect 3384 13880 3390 13932
rect 4522 13880 4528 13932
rect 4580 13920 4586 13932
rect 5123 13923 5181 13929
rect 5123 13920 5135 13923
rect 4580 13892 5135 13920
rect 4580 13880 4586 13892
rect 5123 13889 5135 13892
rect 5169 13920 5181 13923
rect 5442 13920 5448 13932
rect 5169 13892 5448 13920
rect 5169 13889 5181 13892
rect 5123 13883 5181 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 7926 13929 7932 13932
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 5500 13892 6745 13920
rect 5500 13880 5506 13892
rect 6733 13889 6745 13892
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 7920 13883 7932 13929
rect 7926 13880 7932 13883
rect 7984 13880 7990 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10612 13929 10640 13960
rect 10873 13957 10885 13991
rect 10919 13988 10931 13991
rect 11330 13988 11336 14000
rect 10919 13960 11336 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 12406 13960 14320 13988
rect 10778 13929 10784 13932
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10745 13923 10784 13929
rect 10745 13889 10757 13923
rect 10745 13883 10784 13889
rect 1394 13812 1400 13864
rect 1452 13812 1458 13864
rect 1670 13812 1676 13864
rect 1728 13812 1734 13864
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3510 13852 3516 13864
rect 3191 13824 3516 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 3510 13812 3516 13824
rect 3568 13812 3574 13864
rect 3694 13812 3700 13864
rect 3752 13812 3758 13864
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6236 13824 6837 13852
rect 6236 13812 6242 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 7098 13852 7104 13864
rect 6963 13824 7104 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 6932 13784 6960 13815
rect 7098 13812 7104 13824
rect 7156 13812 7162 13864
rect 7650 13812 7656 13864
rect 7708 13812 7714 13864
rect 10042 13812 10048 13864
rect 10100 13812 10106 13864
rect 10612 13852 10640 13883
rect 10778 13880 10784 13883
rect 10836 13880 10842 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 11146 13929 11152 13932
rect 11103 13923 11152 13929
rect 11103 13889 11115 13923
rect 11149 13889 11152 13923
rect 11103 13883 11152 13889
rect 11146 13880 11152 13883
rect 11204 13880 11210 13932
rect 12406 13852 12434 13960
rect 14292 13932 14320 13960
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13920 12679 13923
rect 13262 13920 13268 13932
rect 12667 13892 13268 13920
rect 12667 13889 12679 13892
rect 12621 13883 12679 13889
rect 13262 13880 13268 13892
rect 13320 13920 13326 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13320 13892 14013 13920
rect 13320 13880 13326 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14458 13920 14464 13932
rect 14332 13892 14464 13920
rect 14332 13880 14338 13892
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14642 13929 14648 13932
rect 14609 13923 14648 13929
rect 14609 13889 14621 13923
rect 14609 13883 14648 13889
rect 14642 13880 14648 13883
rect 14700 13880 14706 13932
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 10612 13824 12434 13852
rect 12802 13812 12808 13864
rect 12860 13852 12866 13864
rect 13725 13855 13783 13861
rect 12860 13824 13676 13852
rect 12860 13812 12866 13824
rect 6604 13756 6960 13784
rect 6604 13744 6610 13756
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 11848 13688 12173 13716
rect 11848 13676 11854 13688
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 13648 13716 13676 13824
rect 13725 13821 13737 13855
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13821 13967 13855
rect 14752 13852 14780 13883
rect 14826 13880 14832 13932
rect 14884 13880 14890 13932
rect 14918 13880 14924 13932
rect 14976 13929 14982 13932
rect 14976 13920 14984 13929
rect 15120 13920 15148 14019
rect 17218 14016 17224 14068
rect 17276 14016 17282 14068
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 14976 13892 15021 13920
rect 15120 13892 15945 13920
rect 14976 13883 14984 13892
rect 15933 13889 15945 13892
rect 15979 13889 15991 13923
rect 15933 13883 15991 13889
rect 14976 13880 14982 13883
rect 16114 13880 16120 13932
rect 16172 13880 16178 13932
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 13909 13815 13967 13821
rect 14568 13824 14780 13852
rect 16209 13855 16267 13861
rect 13740 13784 13768 13815
rect 13814 13784 13820 13796
rect 13740 13756 13820 13784
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 13924 13784 13952 13815
rect 14568 13796 14596 13824
rect 16209 13821 16221 13855
rect 16255 13852 16267 13855
rect 17218 13852 17224 13864
rect 16255 13824 17224 13852
rect 16255 13821 16267 13824
rect 16209 13815 16267 13821
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 13998 13784 14004 13796
rect 13924 13756 14004 13784
rect 13998 13744 14004 13756
rect 14056 13744 14062 13796
rect 14550 13744 14556 13796
rect 14608 13744 14614 13796
rect 16298 13784 16304 13796
rect 14660 13756 16304 13784
rect 14660 13716 14688 13756
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 13648 13688 14688 13716
rect 12161 13679 12219 13685
rect 15746 13676 15752 13728
rect 15804 13676 15810 13728
rect 1104 13626 17756 13648
rect 1104 13574 2350 13626
rect 2402 13574 2414 13626
rect 2466 13574 2478 13626
rect 2530 13574 2542 13626
rect 2594 13574 2606 13626
rect 2658 13574 17756 13626
rect 1104 13552 17756 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 1728 13484 2145 13512
rect 1728 13472 1734 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 2133 13475 2191 13481
rect 3694 13472 3700 13524
rect 3752 13512 3758 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3752 13484 3801 13512
rect 3752 13472 3758 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 7926 13472 7932 13524
rect 7984 13472 7990 13524
rect 8294 13472 8300 13524
rect 8352 13472 8358 13524
rect 13262 13472 13268 13524
rect 13320 13472 13326 13524
rect 14921 13515 14979 13521
rect 14921 13481 14933 13515
rect 14967 13512 14979 13515
rect 16022 13512 16028 13524
rect 14967 13484 16028 13512
rect 14967 13481 14979 13484
rect 14921 13475 14979 13481
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 17218 13472 17224 13524
rect 17276 13472 17282 13524
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2188 13348 2697 13376
rect 2188 13336 2194 13348
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 4430 13336 4436 13388
rect 4488 13336 4494 13388
rect 8386 13336 8392 13388
rect 8444 13336 8450 13388
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 9079 13348 11529 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 11517 13345 11529 13348
rect 11563 13376 11575 13379
rect 13262 13376 13268 13388
rect 11563 13348 13268 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 13262 13336 13268 13348
rect 13320 13376 13326 13388
rect 15654 13376 15660 13388
rect 13320 13348 15660 13376
rect 13320 13336 13326 13348
rect 15654 13336 15660 13348
rect 15712 13376 15718 13388
rect 15838 13376 15844 13388
rect 15712 13348 15844 13376
rect 15712 13336 15718 13348
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 3384 13280 5641 13308
rect 3384 13268 3390 13280
rect 5629 13277 5641 13280
rect 5675 13308 5687 13311
rect 5718 13308 5724 13320
rect 5675 13280 5724 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7064 13280 8125 13308
rect 7064 13268 7070 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 14458 13317 14464 13320
rect 14425 13311 14464 13317
rect 14425 13277 14437 13311
rect 14425 13271 14464 13277
rect 14458 13268 14464 13271
rect 14516 13268 14522 13320
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14783 13311 14841 13317
rect 14783 13277 14795 13311
rect 14829 13308 14841 13311
rect 14918 13308 14924 13320
rect 14829 13280 14924 13308
rect 14829 13277 14841 13280
rect 14783 13271 14841 13277
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 16097 13311 16155 13317
rect 16097 13308 16109 13311
rect 15804 13280 16109 13308
rect 15804 13268 15810 13280
rect 16097 13277 16109 13280
rect 16143 13277 16155 13311
rect 16097 13271 16155 13277
rect 2501 13243 2559 13249
rect 2501 13240 2513 13243
rect 1596 13212 2513 13240
rect 1596 13181 1624 13212
rect 2501 13209 2513 13212
rect 2547 13240 2559 13243
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 2547 13212 4169 13240
rect 2547 13209 2559 13212
rect 2501 13203 2559 13209
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 4157 13203 4215 13209
rect 4249 13243 4307 13249
rect 4249 13209 4261 13243
rect 4295 13240 4307 13243
rect 4522 13240 4528 13252
rect 4295 13212 4528 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 7374 13200 7380 13252
rect 7432 13200 7438 13252
rect 9306 13200 9312 13252
rect 9364 13200 9370 13252
rect 10042 13200 10048 13252
rect 10100 13200 10106 13252
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 12526 13200 12532 13252
rect 12584 13200 12590 13252
rect 14642 13200 14648 13252
rect 14700 13200 14706 13252
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 2593 13175 2651 13181
rect 2593 13141 2605 13175
rect 2639 13172 2651 13175
rect 3510 13172 3516 13184
rect 2639 13144 3516 13172
rect 2639 13141 2651 13144
rect 2593 13135 2651 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 10778 13132 10784 13184
rect 10836 13132 10842 13184
rect 1104 13082 17756 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 17756 13082
rect 1104 13008 17756 13030
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 6086 12968 6092 12980
rect 3568 12940 6092 12968
rect 3568 12928 3574 12940
rect 4540 12841 4568 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 7006 12928 7012 12980
rect 7064 12928 7070 12980
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 9364 12940 10057 12968
rect 9364 12928 9370 12940
rect 10045 12937 10057 12940
rect 10091 12937 10103 12971
rect 10045 12931 10103 12937
rect 13262 12928 13268 12980
rect 13320 12928 13326 12980
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 6270 12860 6276 12912
rect 6328 12900 6334 12912
rect 6641 12903 6699 12909
rect 6641 12900 6653 12903
rect 6328 12872 6653 12900
rect 6328 12860 6334 12872
rect 6641 12869 6653 12872
rect 6687 12869 6699 12903
rect 6641 12863 6699 12869
rect 6733 12903 6791 12909
rect 6733 12869 6745 12903
rect 6779 12900 6791 12903
rect 7098 12900 7104 12912
rect 6779 12872 7104 12900
rect 6779 12869 6791 12872
rect 6733 12863 6791 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 17218 12900 17224 12912
rect 16684 12872 17224 12900
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12801 4583 12835
rect 4525 12795 4583 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4663 12804 5764 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4264 12708 4292 12795
rect 4356 12764 4384 12795
rect 5736 12776 5764 12804
rect 5994 12792 6000 12844
rect 6052 12832 6058 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6052 12804 6377 12832
rect 6052 12792 6058 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6454 12792 6460 12844
rect 6512 12792 6518 12844
rect 6822 12792 6828 12844
rect 6880 12841 6886 12844
rect 6880 12835 6907 12841
rect 6895 12801 6907 12835
rect 6880 12795 6907 12801
rect 6880 12792 6886 12795
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10778 12832 10784 12844
rect 10551 12804 10784 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 11790 12792 11796 12844
rect 11848 12792 11854 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13847 12835 13905 12841
rect 13847 12832 13859 12835
rect 13412 12804 13859 12832
rect 13412 12792 13418 12804
rect 13847 12801 13859 12804
rect 13893 12801 13905 12835
rect 13847 12795 13905 12801
rect 13998 12792 14004 12844
rect 14056 12792 14062 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14240 12804 14473 12832
rect 14240 12792 14246 12804
rect 14461 12801 14473 12804
rect 14507 12832 14519 12835
rect 15010 12832 15016 12844
rect 14507 12804 15016 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 16684 12841 16712 12872
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 16669 12835 16727 12841
rect 16669 12801 16681 12835
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 17402 12792 17408 12844
rect 17460 12792 17466 12844
rect 5534 12764 5540 12776
rect 4356 12736 5540 12764
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 10870 12764 10876 12776
rect 10735 12736 10876 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 14918 12764 14924 12776
rect 10928 12736 14924 12764
rect 10928 12724 10934 12736
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 6454 12696 6460 12708
rect 4304 12668 6460 12696
rect 4304 12656 4310 12668
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 13630 12656 13636 12708
rect 13688 12656 13694 12708
rect 13814 12656 13820 12708
rect 13872 12696 13878 12708
rect 17144 12696 17172 12727
rect 13872 12668 17172 12696
rect 13872 12656 13878 12668
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4522 12628 4528 12640
rect 4111 12600 4528 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 14550 12588 14556 12640
rect 14608 12588 14614 12640
rect 16850 12588 16856 12640
rect 16908 12588 16914 12640
rect 1104 12538 17756 12560
rect 1104 12486 2350 12538
rect 2402 12486 2414 12538
rect 2466 12486 2478 12538
rect 2530 12486 2542 12538
rect 2594 12486 2606 12538
rect 2658 12486 17756 12538
rect 1104 12464 17756 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 2924 12396 3157 12424
rect 2924 12384 2930 12396
rect 3145 12393 3157 12396
rect 3191 12424 3203 12427
rect 4246 12424 4252 12436
rect 3191 12396 4252 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 6178 12424 6184 12436
rect 5684 12396 6184 12424
rect 5684 12384 5690 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 7745 12427 7803 12433
rect 7745 12393 7757 12427
rect 7791 12424 7803 12427
rect 7791 12396 7880 12424
rect 7791 12393 7803 12396
rect 7745 12387 7803 12393
rect 7852 12368 7880 12396
rect 12526 12384 12532 12436
rect 12584 12384 12590 12436
rect 15010 12424 15016 12436
rect 14384 12396 15016 12424
rect 4617 12359 4675 12365
rect 4617 12325 4629 12359
rect 4663 12356 4675 12359
rect 5350 12356 5356 12368
rect 4663 12328 5356 12356
rect 4663 12325 4675 12328
rect 4617 12319 4675 12325
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 5810 12356 5816 12368
rect 5592 12328 5816 12356
rect 5592 12316 5598 12328
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 6549 12359 6607 12365
rect 6549 12356 6561 12359
rect 5960 12328 6561 12356
rect 5960 12316 5966 12328
rect 6549 12325 6561 12328
rect 6595 12325 6607 12359
rect 6549 12319 6607 12325
rect 1394 12248 1400 12300
rect 1452 12248 1458 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 4540 12260 6469 12288
rect 3510 12180 3516 12232
rect 3568 12180 3574 12232
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4540 12229 4568 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6564 12288 6592 12319
rect 7834 12316 7840 12368
rect 7892 12316 7898 12368
rect 7926 12316 7932 12368
rect 7984 12316 7990 12368
rect 6564 12260 7834 12288
rect 6457 12251 6515 12257
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4396 12192 4537 12220
rect 4396 12180 4402 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 4890 12220 4896 12232
rect 4847 12192 4896 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 1670 12112 1676 12164
rect 1728 12112 1734 12164
rect 3421 12155 3479 12161
rect 3421 12152 3433 12155
rect 2898 12124 3433 12152
rect 3421 12121 3433 12124
rect 3467 12121 3479 12155
rect 4724 12152 4752 12183
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 5258 12220 5264 12232
rect 5031 12192 5264 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 5534 12220 5540 12232
rect 5495 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12220 5687 12223
rect 5994 12220 6000 12232
rect 5675 12192 6000 12220
rect 5675 12189 5687 12192
rect 5629 12183 5687 12189
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 7190 12220 7196 12232
rect 6963 12192 7196 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7806 12229 7834 12260
rect 7806 12223 7877 12229
rect 7806 12189 7831 12223
rect 7865 12220 7877 12223
rect 8113 12223 8171 12229
rect 7935 12220 8064 12222
rect 8113 12220 8125 12223
rect 7865 12194 8125 12220
rect 7865 12192 7967 12194
rect 8036 12192 8125 12194
rect 7865 12189 7880 12192
rect 7806 12186 7880 12189
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 7819 12183 7877 12186
rect 8113 12183 8171 12189
rect 8202 12180 8208 12232
rect 8260 12180 8266 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 3421 12115 3479 12121
rect 4632 12124 6040 12152
rect 4632 12096 4660 12124
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4341 12087 4399 12093
rect 4341 12084 4353 12087
rect 4304 12056 4353 12084
rect 4304 12044 4310 12056
rect 4341 12053 4353 12056
rect 4387 12053 4399 12087
rect 4341 12047 4399 12053
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5261 12087 5319 12093
rect 5261 12084 5273 12087
rect 5132 12056 5273 12084
rect 5132 12044 5138 12056
rect 5261 12053 5273 12056
rect 5307 12053 5319 12087
rect 5261 12047 5319 12053
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5684 12056 5733 12084
rect 5684 12044 5690 12056
rect 5721 12053 5733 12056
rect 5767 12053 5779 12087
rect 6012 12084 6040 12124
rect 6178 12112 6184 12164
rect 6236 12152 6242 12164
rect 7929 12155 7987 12161
rect 7929 12152 7941 12155
rect 6236 12124 7941 12152
rect 6236 12112 6242 12124
rect 7929 12121 7941 12124
rect 7975 12121 7987 12155
rect 7929 12115 7987 12121
rect 7282 12084 7288 12096
rect 6012 12056 7288 12084
rect 5721 12047 5779 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7834 12084 7840 12096
rect 7524 12056 7840 12084
rect 7524 12044 7530 12056
rect 7834 12044 7840 12056
rect 7892 12084 7898 12096
rect 8312 12084 8340 12183
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 10778 12220 10784 12232
rect 10735 12192 10784 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 14384 12220 14412 12396
rect 15010 12384 15016 12396
rect 15068 12424 15074 12436
rect 15068 12396 16574 12424
rect 15068 12384 15074 12396
rect 16546 12356 16574 12396
rect 16546 12328 16896 12356
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 16669 12291 16727 12297
rect 14516 12260 16528 12288
rect 14516 12248 14522 12260
rect 12483 12192 14412 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 15562 12180 15568 12232
rect 15620 12180 15626 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15896 12192 15945 12220
rect 15896 12180 15902 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 14550 12112 14556 12164
rect 14608 12112 14614 12164
rect 16500 12096 16528 12260
rect 16669 12257 16681 12291
rect 16715 12288 16727 12291
rect 16758 12288 16764 12300
rect 16715 12260 16764 12288
rect 16715 12257 16727 12260
rect 16669 12251 16727 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 16868 12232 16896 12328
rect 16850 12180 16856 12232
rect 16908 12180 16914 12232
rect 7892 12056 8340 12084
rect 7892 12044 7898 12056
rect 8386 12044 8392 12096
rect 8444 12044 8450 12096
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 14139 12087 14197 12093
rect 14139 12053 14151 12087
rect 14185 12084 14197 12087
rect 14734 12084 14740 12096
rect 14185 12056 14740 12084
rect 14185 12053 14197 12056
rect 14139 12047 14197 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15988 12056 16037 12084
rect 15988 12044 15994 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 16390 12044 16396 12096
rect 16448 12044 16454 12096
rect 16482 12044 16488 12096
rect 16540 12044 16546 12096
rect 16942 12044 16948 12096
rect 17000 12044 17006 12096
rect 1104 11994 17756 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 17756 11994
rect 1104 11920 17756 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1728 11852 2145 11880
rect 1728 11840 1734 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 2593 11883 2651 11889
rect 2593 11849 2605 11883
rect 2639 11880 2651 11883
rect 2866 11880 2872 11892
rect 2639 11852 2872 11880
rect 2639 11849 2651 11852
rect 2593 11843 2651 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 5258 11840 5264 11892
rect 5316 11840 5322 11892
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5408 11852 5641 11880
rect 5408 11840 5414 11852
rect 5629 11849 5641 11852
rect 5675 11880 5687 11883
rect 6178 11880 6184 11892
rect 5675 11852 6184 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7340 11852 7757 11880
rect 7340 11840 7346 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 7926 11880 7932 11892
rect 7883 11852 7932 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 13081 11883 13139 11889
rect 13081 11880 13093 11883
rect 12575 11852 13093 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 13081 11849 13093 11852
rect 13127 11849 13139 11883
rect 13081 11843 13139 11849
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 15562 11880 15568 11892
rect 14507 11852 15568 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 2682 11812 2688 11824
rect 2547 11784 2688 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2682 11772 2688 11784
rect 2740 11772 2746 11824
rect 5276 11812 5304 11840
rect 4724 11784 5304 11812
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 4249 11747 4307 11753
rect 2188 11716 2728 11744
rect 2188 11704 2194 11716
rect 2700 11685 2728 11716
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4338 11744 4344 11756
rect 4295 11716 4344 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 4724 11753 4752 11784
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 8113 11815 8171 11821
rect 8113 11812 8125 11815
rect 5592 11784 6224 11812
rect 5592 11772 5598 11784
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5215 11716 5764 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 4614 11676 4620 11688
rect 2685 11639 2743 11645
rect 4356 11648 4620 11676
rect 4356 11617 4384 11648
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 5092 11676 5120 11704
rect 5445 11679 5503 11685
rect 5092 11648 5304 11676
rect 4341 11611 4399 11617
rect 4341 11577 4353 11611
rect 4387 11577 4399 11611
rect 4341 11571 4399 11577
rect 4433 11611 4491 11617
rect 4433 11577 4445 11611
rect 4479 11608 4491 11611
rect 5169 11611 5227 11617
rect 5169 11608 5181 11611
rect 4479 11580 5181 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 5169 11577 5181 11580
rect 5215 11577 5227 11611
rect 5276 11608 5304 11648
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5626 11676 5632 11688
rect 5491 11648 5632 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5736 11676 5764 11716
rect 5810 11704 5816 11756
rect 5868 11704 5874 11756
rect 5920 11753 5948 11784
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 5994 11704 6000 11756
rect 6052 11704 6058 11756
rect 6196 11753 6224 11784
rect 7668 11784 8125 11812
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6454 11744 6460 11756
rect 6227 11716 6460 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 7668 11753 7696 11784
rect 8113 11781 8125 11784
rect 8159 11781 8171 11815
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 8113 11775 8171 11781
rect 8312 11784 12173 11812
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8312 11744 8340 11784
rect 12161 11781 12173 11784
rect 12207 11781 12219 11815
rect 12161 11775 12219 11781
rect 14734 11772 14740 11824
rect 14792 11812 14798 11824
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 14792 11784 14933 11812
rect 14792 11772 14798 11784
rect 14921 11781 14933 11784
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 8067 11716 8340 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 10594 11744 10600 11756
rect 8803 11716 10600 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 5736 11648 6101 11676
rect 6089 11645 6101 11648
rect 6135 11676 6147 11679
rect 8496 11676 8524 11707
rect 6135 11648 8524 11676
rect 6135 11645 6147 11648
rect 6089 11639 6147 11645
rect 8588 11608 8616 11707
rect 10594 11704 10600 11716
rect 10652 11744 10658 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10652 11716 11529 11744
rect 10652 11704 10658 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 11422 11676 11428 11688
rect 8895 11648 11428 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 11422 11636 11428 11648
rect 11480 11676 11486 11688
rect 11624 11676 11652 11707
rect 12066 11704 12072 11756
rect 12124 11704 12130 11756
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12360 11676 12388 11707
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 12710 11704 12716 11756
rect 12768 11744 12774 11756
rect 14752 11744 14780 11772
rect 12768 11716 14780 11744
rect 14829 11747 14887 11753
rect 12768 11704 12774 11716
rect 14829 11713 14841 11747
rect 14875 11744 14887 11747
rect 16114 11744 16120 11756
rect 14875 11716 16120 11744
rect 14875 11713 14887 11716
rect 14829 11707 14887 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17310 11744 17316 11756
rect 17267 11716 17316 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 11480 11648 11652 11676
rect 11900 11648 12388 11676
rect 11480 11636 11486 11648
rect 11900 11617 11928 11648
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12952 11648 13001 11676
rect 12952 11636 12958 11648
rect 12989 11645 13001 11648
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 14182 11676 14188 11688
rect 13127 11648 14188 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14976 11648 15025 11676
rect 14976 11636 14982 11648
rect 15013 11645 15025 11648
rect 15059 11676 15071 11679
rect 16758 11676 16764 11688
rect 15059 11648 16764 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 5276 11580 8616 11608
rect 11885 11611 11943 11617
rect 5169 11571 5227 11577
rect 11885 11577 11897 11611
rect 11931 11577 11943 11611
rect 11885 11571 11943 11577
rect 17402 11568 17408 11620
rect 17460 11568 17466 11620
rect 4062 11500 4068 11552
rect 4120 11500 4126 11552
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 4580 11512 7757 11540
rect 4580 11500 4586 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 11974 11500 11980 11552
rect 12032 11500 12038 11552
rect 12802 11500 12808 11552
rect 12860 11500 12866 11552
rect 1104 11450 17756 11472
rect 1104 11398 2350 11450
rect 2402 11398 2414 11450
rect 2466 11398 2478 11450
rect 2530 11398 2542 11450
rect 2594 11398 2606 11450
rect 2658 11398 17756 11450
rect 1104 11376 17756 11398
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6086 11336 6092 11348
rect 5868 11308 6092 11336
rect 5868 11296 5874 11308
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 10781 11339 10839 11345
rect 10781 11336 10793 11339
rect 7800 11308 10793 11336
rect 7800 11296 7806 11308
rect 10781 11305 10793 11308
rect 10827 11305 10839 11339
rect 10781 11299 10839 11305
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12618 11336 12624 11348
rect 12207 11308 12624 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 12802 11296 12808 11348
rect 12860 11296 12866 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 16540 11308 17417 11336
rect 16540 11296 16546 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 9033 11203 9091 11209
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 11054 11200 11060 11212
rect 9079 11172 11060 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12820 11200 12848 11296
rect 12452 11172 12848 11200
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12452 11141 12480 11172
rect 15930 11160 15936 11212
rect 15988 11160 15994 11212
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12032 11104 12357 11132
rect 12032 11092 12038 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12565 11135 12623 11141
rect 12565 11101 12577 11135
rect 12611 11132 12623 11135
rect 12710 11132 12716 11144
rect 12611 11104 12716 11132
rect 12611 11101 12623 11104
rect 12565 11095 12623 11101
rect 9306 11024 9312 11076
rect 9364 11024 9370 11076
rect 10686 11064 10692 11076
rect 10534 11036 10692 11064
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12161 11067 12219 11073
rect 12161 11064 12173 11067
rect 12124 11036 12173 11064
rect 12124 11024 12130 11036
rect 12161 11033 12173 11036
rect 12207 11064 12219 11067
rect 12360 11064 12388 11095
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12860 11104 12909 11132
rect 12860 11092 12866 11104
rect 12897 11101 12909 11104
rect 12943 11132 12955 11135
rect 13722 11132 13728 11144
rect 12943 11104 13728 11132
rect 12943 11101 12955 11104
rect 12897 11095 12955 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 15620 11104 15669 11132
rect 15620 11092 15626 11104
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 14458 11064 14464 11076
rect 12207 11036 12296 11064
rect 12360 11036 14464 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 1581 10999 1639 11005
rect 1581 10965 1593 10999
rect 1627 10996 1639 10999
rect 2682 10996 2688 11008
rect 1627 10968 2688 10996
rect 1627 10965 1639 10968
rect 1581 10959 1639 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 9030 10996 9036 11008
rect 4580 10968 9036 10996
rect 4580 10956 4586 10968
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 12268 10996 12296 11036
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 16942 11024 16948 11076
rect 17000 11024 17006 11076
rect 12434 10996 12440 11008
rect 12268 10968 12440 10996
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 17756 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 17756 10906
rect 1104 10832 17756 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2682 10792 2688 10804
rect 2547 10764 2688 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5718 10752 5724 10804
rect 5776 10752 5782 10804
rect 7098 10752 7104 10804
rect 7156 10752 7162 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 7432 10764 10057 10792
rect 7432 10752 7438 10764
rect 10045 10761 10057 10764
rect 10091 10792 10103 10795
rect 11790 10792 11796 10804
rect 10091 10764 11796 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 13630 10792 13636 10804
rect 13219 10764 13636 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14826 10792 14832 10804
rect 14599 10764 14832 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 17221 10795 17279 10801
rect 17221 10792 17233 10795
rect 16172 10764 17233 10792
rect 16172 10752 16178 10764
rect 17221 10761 17233 10764
rect 17267 10761 17279 10795
rect 17221 10755 17279 10761
rect 1302 10684 1308 10736
rect 1360 10724 1366 10736
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 1360 10696 8769 10724
rect 1360 10684 1366 10696
rect 8757 10693 8769 10696
rect 8803 10693 8815 10727
rect 8757 10687 8815 10693
rect 10686 10684 10692 10736
rect 10744 10684 10750 10736
rect 13648 10696 14320 10724
rect 2593 10659 2651 10665
rect 2593 10625 2605 10659
rect 2639 10656 2651 10659
rect 3142 10656 3148 10668
rect 2639 10628 3148 10656
rect 2639 10625 2651 10628
rect 2593 10619 2651 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2685 10591 2743 10597
rect 2685 10588 2697 10591
rect 2280 10560 2697 10588
rect 2280 10548 2286 10560
rect 2685 10557 2697 10560
rect 2731 10557 2743 10591
rect 4172 10588 4200 10619
rect 4246 10616 4252 10668
rect 4304 10616 4310 10668
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10656 4399 10659
rect 4430 10656 4436 10668
rect 4387 10628 4436 10656
rect 4387 10625 4399 10628
rect 4341 10619 4399 10625
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 4847 10628 5304 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4172 10560 4629 10588
rect 2685 10551 2743 10557
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 4985 10591 5043 10597
rect 4985 10557 4997 10591
rect 5031 10557 5043 10591
rect 5276 10588 5304 10628
rect 5350 10616 5356 10668
rect 5408 10665 5414 10668
rect 5408 10659 5441 10665
rect 5429 10625 5441 10659
rect 5408 10619 5441 10625
rect 5408 10616 5414 10619
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 5960 10628 6745 10656
rect 5960 10616 5966 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6972 10628 7205 10656
rect 6972 10616 6978 10628
rect 5552 10588 5580 10616
rect 5276 10560 5580 10588
rect 4985 10551 5043 10557
rect 5000 10520 5028 10551
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 5534 10520 5540 10532
rect 5000 10492 5540 10520
rect 5534 10480 5540 10492
rect 5592 10520 5598 10532
rect 5994 10520 6000 10532
rect 5592 10492 6000 10520
rect 5592 10480 5598 10492
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 1670 10412 1676 10464
rect 1728 10452 1734 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 1728 10424 2145 10452
rect 1728 10412 1734 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 3881 10455 3939 10461
rect 3881 10452 3893 10455
rect 3568 10424 3893 10452
rect 3568 10412 3574 10424
rect 3881 10421 3893 10424
rect 3927 10421 3939 10455
rect 3881 10415 3939 10421
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 5350 10452 5356 10464
rect 4028 10424 5356 10452
rect 4028 10412 4034 10424
rect 5350 10412 5356 10424
rect 5408 10452 5414 10464
rect 6656 10452 6684 10551
rect 5408 10424 6684 10452
rect 7116 10452 7144 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7331 10628 7696 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 7668 10588 7696 10628
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7834 10616 7840 10668
rect 7892 10616 7898 10668
rect 9950 10616 9956 10668
rect 10008 10656 10014 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 10008 10628 10793 10656
rect 10008 10616 10014 10628
rect 10781 10625 10793 10628
rect 10827 10656 10839 10659
rect 10870 10656 10876 10668
rect 10827 10628 10876 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 13648 10665 13676 10696
rect 11977 10659 12035 10665
rect 11977 10656 11989 10659
rect 11296 10628 11989 10656
rect 11296 10616 11302 10628
rect 11977 10625 11989 10628
rect 12023 10656 12035 10659
rect 12989 10659 13047 10665
rect 12023 10628 12434 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 7852 10588 7880 10616
rect 7668 10560 7880 10588
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 7377 10523 7435 10529
rect 7377 10520 7389 10523
rect 7248 10492 7389 10520
rect 7248 10480 7254 10492
rect 7377 10489 7389 10492
rect 7423 10489 7435 10523
rect 7377 10483 7435 10489
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 8110 10520 8116 10532
rect 7800 10492 8116 10520
rect 7800 10480 7806 10492
rect 8110 10480 8116 10492
rect 8168 10480 8174 10532
rect 12406 10520 12434 10628
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 13357 10659 13415 10665
rect 13357 10656 13369 10659
rect 13311 10628 13369 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 13357 10625 13369 10628
rect 13403 10625 13415 10659
rect 13357 10619 13415 10625
rect 13632 10659 13690 10665
rect 13632 10625 13644 10659
rect 13678 10625 13690 10659
rect 13632 10619 13690 10625
rect 13004 10588 13032 10619
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 14292 10665 14320 10696
rect 14277 10659 14335 10665
rect 13780 10628 13952 10656
rect 13780 10616 13786 10628
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 13004 10560 13829 10588
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 13924 10588 13952 10628
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14323 10628 14933 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 14967 10628 16252 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 16224 10600 16252 10628
rect 17126 10616 17132 10668
rect 17184 10616 17190 10668
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 13924 10560 15025 10588
rect 13924 10529 13952 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 16206 10548 16212 10600
rect 16264 10548 16270 10600
rect 16298 10548 16304 10600
rect 16356 10548 16362 10600
rect 13909 10523 13967 10529
rect 12406 10492 13124 10520
rect 8294 10452 8300 10464
rect 7116 10424 8300 10452
rect 5408 10412 5414 10424
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 12032 10424 12081 10452
rect 12032 10412 12038 10424
rect 12069 10421 12081 10424
rect 12115 10452 12127 10455
rect 12894 10452 12900 10464
rect 12115 10424 12900 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 12986 10412 12992 10464
rect 13044 10412 13050 10464
rect 13096 10452 13124 10492
rect 13909 10489 13921 10523
rect 13955 10489 13967 10523
rect 16945 10523 17003 10529
rect 16945 10520 16957 10523
rect 13909 10483 13967 10489
rect 15120 10492 16957 10520
rect 15120 10464 15148 10492
rect 16945 10489 16957 10492
rect 16991 10489 17003 10523
rect 16945 10483 17003 10489
rect 13998 10452 14004 10464
rect 13096 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 15102 10412 15108 10464
rect 15160 10412 15166 10464
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 15838 10452 15844 10464
rect 15795 10424 15844 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 1104 10362 17756 10384
rect 1104 10310 2350 10362
rect 2402 10310 2414 10362
rect 2466 10310 2478 10362
rect 2530 10310 2542 10362
rect 2594 10310 2606 10362
rect 2658 10310 17756 10362
rect 1104 10288 17756 10310
rect 5261 10251 5319 10257
rect 5261 10217 5273 10251
rect 5307 10248 5319 10251
rect 5534 10248 5540 10260
rect 5307 10220 5540 10248
rect 5307 10217 5319 10220
rect 5261 10211 5319 10217
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7742 10248 7748 10260
rect 7524 10220 7748 10248
rect 7524 10208 7530 10220
rect 7742 10208 7748 10220
rect 7800 10248 7806 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 7800 10220 8309 10248
rect 7800 10208 7806 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 10962 10208 10968 10260
rect 11020 10208 11026 10260
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 16264 10220 17325 10248
rect 16264 10208 16270 10220
rect 17313 10217 17325 10220
rect 17359 10217 17371 10251
rect 17313 10211 17371 10217
rect 3786 10140 3792 10192
rect 3844 10140 3850 10192
rect 4080 10152 6132 10180
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 2866 10112 2872 10124
rect 1443 10084 2872 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2866 10072 2872 10084
rect 2924 10112 2930 10124
rect 4080 10112 4108 10152
rect 5902 10112 5908 10124
rect 2924 10084 4108 10112
rect 5276 10084 5908 10112
rect 2924 10072 2930 10084
rect 3418 10004 3424 10056
rect 3476 10004 3482 10056
rect 4062 10004 4068 10056
rect 4120 10004 4126 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4522 10044 4528 10056
rect 4479 10016 4528 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4522 10004 4528 10016
rect 4580 10044 4586 10056
rect 5074 10044 5080 10056
rect 4580 10016 5080 10044
rect 4580 10004 4586 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5186 10047 5244 10053
rect 5186 10013 5198 10047
rect 5232 10044 5244 10047
rect 5276 10044 5304 10084
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 5232 10016 5304 10044
rect 5232 10013 5244 10016
rect 5186 10007 5244 10013
rect 5442 10004 5448 10056
rect 5500 10004 5506 10056
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5718 10044 5724 10056
rect 5583 10016 5724 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6104 10053 6132 10152
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7558 10112 7564 10124
rect 7340 10084 7564 10112
rect 7340 10072 7346 10084
rect 7558 10072 7564 10084
rect 7616 10112 7622 10124
rect 7616 10084 8248 10112
rect 7616 10072 7622 10084
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6914 10044 6920 10056
rect 6135 10016 6920 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8220 10053 8248 10084
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11422 10112 11428 10124
rect 11020 10084 11428 10112
rect 11020 10072 11026 10084
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 13814 10112 13820 10124
rect 11655 10084 13820 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 13814 10072 13820 10084
rect 13872 10112 13878 10124
rect 15010 10112 15016 10124
rect 13872 10084 15016 10112
rect 13872 10072 13878 10084
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15838 10072 15844 10124
rect 15896 10072 15902 10124
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 8076 10016 8125 10044
rect 8076 10004 8082 10016
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8206 10047 8264 10053
rect 8206 10013 8218 10047
rect 8252 10013 8264 10047
rect 8206 10007 8264 10013
rect 11790 10004 11796 10056
rect 11848 10004 11854 10056
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 1670 9936 1676 9988
rect 1728 9936 1734 9988
rect 3329 9979 3387 9985
rect 3329 9976 3341 9979
rect 2898 9948 3341 9976
rect 3329 9945 3341 9948
rect 3375 9945 3387 9979
rect 3329 9939 3387 9945
rect 3789 9979 3847 9985
rect 3789 9945 3801 9979
rect 3835 9976 3847 9979
rect 4341 9979 4399 9985
rect 4341 9976 4353 9979
rect 3835 9948 4353 9976
rect 3835 9945 3847 9948
rect 3789 9939 3847 9945
rect 4341 9945 4353 9948
rect 4387 9976 4399 9979
rect 9122 9976 9128 9988
rect 4387 9948 9128 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 16574 9936 16580 9988
rect 16632 9936 16638 9988
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3878 9908 3884 9920
rect 3200 9880 3884 9908
rect 3200 9868 3206 9880
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 3973 9911 4031 9917
rect 3973 9877 3985 9911
rect 4019 9908 4031 9911
rect 4430 9908 4436 9920
rect 4019 9880 4436 9908
rect 4019 9877 4031 9880
rect 3973 9871 4031 9877
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 5684 9880 5733 9908
rect 5684 9868 5690 9880
rect 5721 9877 5733 9880
rect 5767 9877 5779 9911
rect 5721 9871 5779 9877
rect 11330 9868 11336 9920
rect 11388 9868 11394 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 13081 9911 13139 9917
rect 13081 9908 13093 9911
rect 11848 9880 13093 9908
rect 11848 9868 11854 9880
rect 13081 9877 13093 9880
rect 13127 9877 13139 9911
rect 13081 9871 13139 9877
rect 1104 9818 17756 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 17756 9818
rect 1104 9744 17756 9766
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 5902 9704 5908 9716
rect 3936 9676 5908 9704
rect 3936 9664 3942 9676
rect 5902 9664 5908 9676
rect 5960 9664 5966 9716
rect 6825 9707 6883 9713
rect 6825 9673 6837 9707
rect 6871 9704 6883 9707
rect 6914 9704 6920 9716
rect 6871 9676 6920 9704
rect 6871 9673 6883 9676
rect 6825 9667 6883 9673
rect 6914 9664 6920 9676
rect 6972 9704 6978 9716
rect 7650 9704 7656 9716
rect 6972 9676 7656 9704
rect 6972 9664 6978 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 7432 9608 8125 9636
rect 7432 9596 7438 9608
rect 8113 9605 8125 9608
rect 8159 9605 8171 9639
rect 8113 9599 8171 9605
rect 9306 9596 9312 9648
rect 9364 9636 9370 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 9364 9608 9505 9636
rect 9364 9596 9370 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9769 9639 9827 9645
rect 9769 9605 9781 9639
rect 9815 9636 9827 9639
rect 11072 9636 11100 9667
rect 9815 9608 10180 9636
rect 11072 9608 11928 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 10152 9580 10180 9608
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9232 9540 9597 9568
rect 9232 9512 9260 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9916 9540 9965 9568
rect 9916 9528 9922 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 9953 9531 10011 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10597 9571 10655 9577
rect 10597 9568 10609 9571
rect 10459 9540 10609 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10597 9537 10609 9540
rect 10643 9537 10655 9571
rect 10597 9531 10655 9537
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 10962 9568 10968 9580
rect 10919 9540 10968 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11790 9568 11796 9580
rect 11112 9540 11796 9568
rect 11112 9528 11118 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 11900 9568 11928 9608
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 13449 9639 13507 9645
rect 13449 9636 13461 9639
rect 12492 9608 13461 9636
rect 12492 9596 12498 9608
rect 13449 9605 13461 9608
rect 13495 9605 13507 9639
rect 13449 9599 13507 9605
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16632 9608 16773 9636
rect 16632 9596 16638 9608
rect 16761 9605 16773 9608
rect 16807 9605 16819 9639
rect 16761 9599 16819 9605
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 11900 9540 13553 9568
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 14783 9540 16574 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9048 9364 9076 9463
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 10321 9503 10379 9509
rect 10321 9500 10333 9503
rect 9355 9472 10333 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 10321 9469 10333 9472
rect 10367 9469 10379 9503
rect 10321 9463 10379 9469
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 9582 9392 9588 9444
rect 9640 9392 9646 9444
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 9048 9336 10057 9364
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 11164 9364 11192 9463
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 11480 9472 12817 9500
rect 11480 9460 11486 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 13556 9500 13584 9531
rect 13906 9500 13912 9512
rect 13556 9472 13912 9500
rect 12805 9463 12863 9469
rect 13906 9460 13912 9472
rect 13964 9500 13970 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 13964 9472 14841 9500
rect 13964 9460 13970 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 15010 9460 15016 9512
rect 15068 9460 15074 9512
rect 16546 9500 16574 9540
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 16758 9500 16764 9512
rect 16546 9472 16764 9500
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 11330 9392 11336 9444
rect 11388 9432 11394 9444
rect 13173 9435 13231 9441
rect 13173 9432 13185 9435
rect 11388 9404 13185 9432
rect 11388 9392 11394 9404
rect 13173 9401 13185 9404
rect 13219 9432 13231 9435
rect 13538 9432 13544 9444
rect 13219 9404 13544 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 14369 9435 14427 9441
rect 14369 9401 14381 9435
rect 14415 9432 14427 9435
rect 14642 9432 14648 9444
rect 14415 9404 14648 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 17221 9435 17279 9441
rect 17221 9432 17233 9435
rect 16448 9404 17233 9432
rect 16448 9392 16454 9404
rect 17221 9401 17233 9404
rect 17267 9401 17279 9435
rect 17221 9395 17279 9401
rect 12526 9364 12532 9376
rect 11164 9336 12532 9364
rect 10045 9327 10103 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 12768 9336 13277 9364
rect 12768 9324 12774 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 1104 9274 17756 9296
rect 1104 9222 2350 9274
rect 2402 9222 2414 9274
rect 2466 9222 2478 9274
rect 2530 9222 2542 9274
rect 2594 9222 2606 9274
rect 2658 9222 17756 9274
rect 1104 9200 17756 9222
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 9214 9160 9220 9172
rect 5859 9132 9220 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 10226 9160 10232 9172
rect 9364 9132 10232 9160
rect 9364 9120 9370 9132
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13044 9132 13369 9160
rect 13044 9120 13050 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 3970 9052 3976 9104
rect 4028 9052 4034 9104
rect 7285 9095 7343 9101
rect 7285 9061 7297 9095
rect 7331 9092 7343 9095
rect 9858 9092 9864 9104
rect 7331 9064 9864 9092
rect 7331 9061 7343 9064
rect 7285 9055 7343 9061
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 12710 9052 12716 9104
rect 12768 9052 12774 9104
rect 13998 9092 14004 9104
rect 13004 9064 14004 9092
rect 3878 8916 3884 8968
rect 3936 8916 3942 8968
rect 3988 8965 4016 9052
rect 5718 8984 5724 9036
rect 5776 8984 5782 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6638 9024 6644 9036
rect 5859 8996 6644 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6638 8984 6644 8996
rect 6696 9024 6702 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6696 8996 6929 9024
rect 6696 8984 6702 8996
rect 6917 8993 6929 8996
rect 6963 8993 6975 9027
rect 7466 9024 7472 9036
rect 6917 8987 6975 8993
rect 7024 8996 7472 9024
rect 3974 8959 4032 8965
rect 3974 8925 3986 8959
rect 4020 8925 4032 8959
rect 3974 8919 4032 8925
rect 3878 8780 3884 8832
rect 3936 8820 3942 8832
rect 3988 8820 4016 8919
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 7024 8965 7052 8996
rect 7466 8984 7472 8996
rect 7524 9024 7530 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7524 8996 7573 9024
rect 7524 8984 7530 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 7742 9024 7748 9036
rect 7699 8996 7748 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 7834 8984 7840 9036
rect 7892 9024 7898 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7892 8996 8033 9024
rect 7892 8984 7898 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 10778 9024 10784 9036
rect 8021 8987 8079 8993
rect 8220 8996 10784 9024
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 5997 8891 6055 8897
rect 5997 8888 6009 8891
rect 4856 8860 6009 8888
rect 4856 8848 4862 8860
rect 5997 8857 6009 8860
rect 6043 8857 6055 8891
rect 6840 8888 6868 8919
rect 7098 8916 7104 8968
rect 7156 8916 7162 8968
rect 7190 8916 7196 8968
rect 7248 8916 7254 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 7208 8888 7236 8916
rect 6840 8860 7236 8888
rect 7300 8888 7328 8919
rect 7469 8891 7527 8897
rect 7469 8888 7481 8891
rect 7300 8860 7481 8888
rect 5997 8851 6055 8857
rect 7469 8857 7481 8860
rect 7515 8857 7527 8891
rect 7944 8888 7972 8919
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8220 8965 8248 8996
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8168 8928 8217 8956
rect 8168 8916 8174 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8680 8965 8708 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12805 9027 12863 9033
rect 12805 9024 12817 9027
rect 12492 8996 12817 9024
rect 12492 8984 12498 8996
rect 12805 8993 12817 8996
rect 12851 8993 12863 9027
rect 12805 8987 12863 8993
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8352 8928 8493 8956
rect 8352 8916 8358 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13004 8956 13032 9064
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 13173 9027 13231 9033
rect 13173 8993 13185 9027
rect 13219 9024 13231 9027
rect 15381 9027 15439 9033
rect 13219 8996 13308 9024
rect 13219 8993 13231 8996
rect 13173 8987 13231 8993
rect 12943 8928 13032 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 8018 8888 8024 8900
rect 7944 8860 8024 8888
rect 7469 8851 7527 8857
rect 3936 8792 4016 8820
rect 4249 8823 4307 8829
rect 3936 8780 3942 8792
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 4522 8820 4528 8832
rect 4295 8792 4528 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 6012 8820 6040 8851
rect 8018 8848 8024 8860
rect 8076 8888 8082 8900
rect 8573 8891 8631 8897
rect 8573 8888 8585 8891
rect 8076 8860 8585 8888
rect 8076 8848 8082 8860
rect 8573 8857 8585 8860
rect 8619 8857 8631 8891
rect 8573 8851 8631 8857
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 10192 8860 13185 8888
rect 10192 8848 10198 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 7006 8820 7012 8832
rect 6012 8792 7012 8820
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13081 8823 13139 8829
rect 13081 8820 13093 8823
rect 12860 8792 13093 8820
rect 12860 8780 12866 8792
rect 13081 8789 13093 8792
rect 13127 8820 13139 8823
rect 13280 8820 13308 8996
rect 15381 8993 15393 9027
rect 15427 9024 15439 9027
rect 16298 9024 16304 9036
rect 15427 8996 16304 9024
rect 15427 8993 15439 8996
rect 15381 8987 15439 8993
rect 16298 8984 16304 8996
rect 16356 9024 16362 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16356 8996 16589 9024
rect 16356 8984 16362 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 13446 8916 13452 8968
rect 13504 8916 13510 8968
rect 15102 8916 15108 8968
rect 15160 8916 15166 8968
rect 16390 8916 16396 8968
rect 16448 8916 16454 8968
rect 13538 8848 13544 8900
rect 13596 8888 13602 8900
rect 13596 8860 15240 8888
rect 13596 8848 13602 8860
rect 13127 8792 13308 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 15212 8829 15240 8860
rect 14737 8823 14795 8829
rect 14737 8820 14749 8823
rect 14608 8792 14749 8820
rect 14608 8780 14614 8792
rect 14737 8789 14749 8792
rect 14783 8789 14795 8823
rect 14737 8783 14795 8789
rect 15197 8823 15255 8829
rect 15197 8789 15209 8823
rect 15243 8820 15255 8823
rect 15838 8820 15844 8832
rect 15243 8792 15844 8820
rect 15243 8789 15255 8792
rect 15197 8783 15255 8789
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15988 8792 16037 8820
rect 15988 8780 15994 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16758 8820 16764 8832
rect 16531 8792 16764 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 1104 8730 17756 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 17756 8730
rect 1104 8656 17756 8678
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 2608 8588 3341 8616
rect 2608 8548 2636 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 3528 8588 5396 8616
rect 2438 8520 2636 8548
rect 2866 8508 2872 8560
rect 2924 8548 2930 8560
rect 2924 8520 3188 8548
rect 2924 8508 2930 8520
rect 3160 8489 3188 8520
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3528 8480 3556 8588
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 3651 8520 4108 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 4080 8489 4108 8520
rect 3819 8483 3877 8489
rect 3819 8480 3831 8483
rect 3528 8452 3831 8480
rect 3819 8449 3831 8452
rect 3865 8449 3877 8483
rect 3819 8443 3877 8449
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3510 8412 3516 8424
rect 2915 8384 3516 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3510 8372 3516 8384
rect 3568 8372 3574 8424
rect 3988 8344 4016 8443
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4522 8440 4528 8492
rect 4580 8440 4586 8492
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5368 8489 5396 8588
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5776 8588 6009 8616
rect 5776 8576 5782 8588
rect 5997 8585 6009 8588
rect 6043 8585 6055 8619
rect 5997 8579 6055 8585
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4939 8452 4997 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5260 8483 5318 8489
rect 5260 8449 5272 8483
rect 5306 8449 5318 8483
rect 5260 8443 5318 8449
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5442 8480 5448 8492
rect 5399 8452 5448 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5276 8344 5304 8443
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5902 8480 5908 8492
rect 5859 8452 5908 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6012 8480 6040 8579
rect 7926 8576 7932 8628
rect 7984 8576 7990 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12618 8616 12624 8628
rect 11931 8588 12624 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12618 8576 12624 8588
rect 12676 8616 12682 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 12676 8588 13369 8616
rect 12676 8576 12682 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 7944 8548 7972 8576
rect 7392 8520 7972 8548
rect 6012 8452 6500 8480
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5592 8384 5641 8412
rect 5592 8372 5598 8384
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 6472 8421 6500 8452
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7006 8480 7012 8492
rect 6779 8452 7012 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7392 8489 7420 8520
rect 7668 8489 7696 8520
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 13449 8551 13507 8557
rect 11480 8520 11652 8548
rect 11480 8508 11486 8520
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5776 8384 6377 8412
rect 5776 8372 5782 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 6457 8415 6515 8421
rect 6457 8381 6469 8415
rect 6503 8381 6515 8415
rect 7576 8412 7604 8443
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7892 8452 7941 8480
rect 7892 8440 7898 8452
rect 7929 8449 7941 8452
rect 7975 8449 7987 8483
rect 7929 8443 7987 8449
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 11624 8489 11652 8520
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13633 8551 13691 8557
rect 13633 8548 13645 8551
rect 13495 8520 13645 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13633 8517 13645 8520
rect 13679 8517 13691 8551
rect 13633 8511 13691 8517
rect 13924 8520 14596 8548
rect 13924 8492 13952 8520
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11388 8452 11529 8480
rect 11388 8440 11394 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11610 8483 11668 8489
rect 11610 8449 11622 8483
rect 11656 8449 11668 8483
rect 11610 8443 11668 8449
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13906 8480 13912 8492
rect 13867 8452 13912 8480
rect 13541 8443 13599 8449
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7576 8384 7757 8412
rect 6457 8375 6515 8381
rect 7745 8381 7757 8384
rect 7791 8412 7803 8415
rect 8202 8412 8208 8424
rect 7791 8384 8208 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 5810 8344 5816 8356
rect 3988 8316 5816 8344
rect 5810 8304 5816 8316
rect 5868 8344 5874 8356
rect 6546 8344 6552 8356
rect 5868 8316 6552 8344
rect 5868 8304 5874 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 6880 8316 6929 8344
rect 6880 8304 6886 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 12618 8304 12624 8356
rect 12676 8304 12682 8356
rect 13096 8344 13124 8443
rect 13170 8372 13176 8424
rect 13228 8372 13234 8424
rect 13556 8412 13584 8443
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14568 8489 14596 8520
rect 14460 8483 14518 8489
rect 14460 8480 14472 8483
rect 14056 8452 14472 8480
rect 14056 8440 14062 8452
rect 14460 8449 14472 8452
rect 14506 8449 14518 8483
rect 14460 8443 14518 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13556 8384 14197 8412
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14476 8412 14504 8443
rect 16758 8412 16764 8424
rect 14476 8384 16764 8412
rect 14185 8375 14243 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 13446 8344 13452 8356
rect 13096 8316 13452 8344
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 1397 8279 1455 8285
rect 1397 8245 1409 8279
rect 1443 8276 1455 8279
rect 1578 8276 1584 8288
rect 1443 8248 1584 8276
rect 1443 8245 1455 8248
rect 1397 8239 1455 8245
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 7466 8236 7472 8288
rect 7524 8236 7530 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 8076 8248 8217 8276
rect 8076 8236 8082 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 1104 8186 17756 8208
rect 1104 8134 2350 8186
rect 2402 8134 2414 8186
rect 2466 8134 2478 8186
rect 2530 8134 2542 8186
rect 2594 8134 2606 8186
rect 2658 8134 17756 8186
rect 1104 8112 17756 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 1397 8075 1455 8081
rect 1397 8072 1409 8075
rect 1360 8044 1409 8072
rect 1360 8032 1366 8044
rect 1397 8041 1409 8044
rect 1443 8041 1455 8075
rect 1397 8035 1455 8041
rect 12253 8075 12311 8081
rect 12253 8041 12265 8075
rect 12299 8072 12311 8075
rect 13170 8072 13176 8084
rect 12299 8044 13176 8072
rect 12299 8041 12311 8044
rect 12253 8035 12311 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 17359 8075 17417 8081
rect 17359 8072 17371 8075
rect 16816 8044 17371 8072
rect 16816 8032 16822 8044
rect 17359 8041 17371 8044
rect 17405 8041 17417 8075
rect 17359 8035 17417 8041
rect 4246 7964 4252 8016
rect 4304 7964 4310 8016
rect 10689 8007 10747 8013
rect 10689 7973 10701 8007
rect 10735 8004 10747 8007
rect 12618 8004 12624 8016
rect 10735 7976 12624 8004
rect 10735 7973 10747 7976
rect 10689 7967 10747 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 7156 7908 10793 7936
rect 7156 7896 7162 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11388 7908 12204 7936
rect 11388 7896 11394 7908
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 3878 7828 3884 7880
rect 3936 7828 3942 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 6917 7871 6975 7877
rect 4028 7840 4073 7868
rect 4028 7828 4034 7840
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7006 7868 7012 7880
rect 6963 7840 7012 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 8018 7828 8024 7880
rect 8076 7828 8082 7880
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10284 7840 10333 7868
rect 10284 7828 10290 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 12176 7877 12204 7908
rect 15930 7896 15936 7948
rect 15988 7896 15994 7948
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11480 7840 12081 7868
rect 11480 7828 11486 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12162 7871 12220 7877
rect 12162 7837 12174 7871
rect 12208 7837 12220 7871
rect 12162 7831 12220 7837
rect 15562 7828 15568 7880
rect 15620 7828 15626 7880
rect 10505 7803 10563 7809
rect 10505 7769 10517 7803
rect 10551 7800 10563 7803
rect 11974 7800 11980 7812
rect 10551 7772 11980 7800
rect 10551 7769 10563 7772
rect 10505 7763 10563 7769
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 16758 7760 16764 7812
rect 16816 7760 16822 7812
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1673 7735 1731 7741
rect 1673 7732 1685 7735
rect 900 7704 1685 7732
rect 900 7692 906 7704
rect 1673 7701 1685 7704
rect 1719 7701 1731 7735
rect 1673 7695 1731 7701
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 9640 7704 10057 7732
rect 9640 7692 9646 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10413 7735 10471 7741
rect 10413 7701 10425 7735
rect 10459 7732 10471 7735
rect 10778 7732 10784 7744
rect 10459 7704 10784 7732
rect 10459 7701 10471 7704
rect 10413 7695 10471 7701
rect 10778 7692 10784 7704
rect 10836 7692 10842 7744
rect 1104 7642 17756 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 17756 7642
rect 1104 7568 17756 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 1854 7528 1860 7540
rect 1443 7500 1860 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 11054 7528 11060 7540
rect 9416 7500 11060 7528
rect 2222 7420 2228 7472
rect 2280 7420 2286 7472
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 8128 7460 8156 7488
rect 9416 7460 9444 7500
rect 11054 7488 11060 7500
rect 11112 7528 11118 7540
rect 12434 7528 12440 7540
rect 11112 7500 12440 7528
rect 11112 7488 11118 7500
rect 12434 7488 12440 7500
rect 12492 7528 12498 7540
rect 15562 7528 15568 7540
rect 12492 7500 15568 7528
rect 12492 7488 12498 7500
rect 2924 7432 3188 7460
rect 8128 7432 9168 7460
rect 2924 7420 2930 7432
rect 3160 7401 3188 7432
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 4890 7392 4896 7404
rect 3191 7364 4896 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 9140 7401 9168 7432
rect 9324 7432 9444 7460
rect 9324 7401 9352 7432
rect 9582 7420 9588 7472
rect 9640 7420 9646 7472
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 11333 7463 11391 7469
rect 11333 7460 11345 7463
rect 11296 7432 11345 7460
rect 11296 7420 11302 7432
rect 11333 7429 11345 7432
rect 11379 7429 11391 7463
rect 11333 7423 11391 7429
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7524 7364 8125 7392
rect 7524 7352 7530 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3786 7324 3792 7336
rect 2915 7296 3792 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 9048 7324 9076 7355
rect 10686 7352 10692 7404
rect 10744 7352 10750 7404
rect 14292 7401 14320 7500
rect 15562 7488 15568 7500
rect 15620 7488 15626 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15896 7500 16037 7528
rect 15896 7488 15902 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 16758 7488 16764 7540
rect 16816 7488 16822 7540
rect 14550 7420 14556 7472
rect 14608 7420 14614 7472
rect 16209 7463 16267 7469
rect 16209 7460 16221 7463
rect 15778 7432 16221 7460
rect 16209 7429 16221 7432
rect 16255 7429 16267 7463
rect 16209 7423 16267 7429
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16850 7392 16856 7404
rect 16347 7364 16381 7392
rect 16546 7364 16856 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 9582 7324 9588 7336
rect 9048 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7324 9646 7336
rect 11422 7324 11428 7336
rect 9640 7296 11428 7324
rect 9640 7284 9646 7296
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 16316 7324 16344 7355
rect 16546 7324 16574 7364
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 15252 7296 16574 7324
rect 15252 7284 15258 7296
rect 8849 7191 8907 7197
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 8938 7188 8944 7200
rect 8895 7160 8944 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 1104 7098 17756 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 17756 7098
rect 1104 7024 17756 7046
rect 8202 6944 8208 6996
rect 8260 6944 8266 6996
rect 5626 6916 5632 6928
rect 5460 6888 5632 6916
rect 2222 6808 2228 6860
rect 2280 6848 2286 6860
rect 2593 6851 2651 6857
rect 2593 6848 2605 6851
rect 2280 6820 2605 6848
rect 2280 6808 2286 6820
rect 2593 6817 2605 6820
rect 2639 6817 2651 6851
rect 2593 6811 2651 6817
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 5460 6848 5488 6888
rect 5626 6876 5632 6888
rect 5684 6876 5690 6928
rect 8220 6916 8248 6944
rect 8220 6888 8340 6916
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 4479 6820 5488 6848
rect 5552 6820 5733 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 3418 6780 3424 6792
rect 2731 6752 3424 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 3418 6740 3424 6752
rect 3476 6780 3482 6792
rect 3786 6780 3792 6792
rect 3476 6752 3792 6780
rect 3476 6740 3482 6752
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3936 6752 4353 6780
rect 3936 6740 3942 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 4356 6644 4384 6743
rect 5368 6712 5396 6743
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5552 6789 5580 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8202 6848 8208 6860
rect 8159 6820 8208 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 5537 6783 5595 6789
rect 5537 6749 5549 6783
rect 5583 6749 5595 6783
rect 5537 6743 5595 6749
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6089 6715 6147 6721
rect 6089 6712 6101 6715
rect 5368 6684 6101 6712
rect 6089 6681 6101 6684
rect 6135 6681 6147 6715
rect 6089 6675 6147 6681
rect 6196 6644 6224 6743
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 6604 6752 6653 6780
rect 6604 6740 6610 6752
rect 6641 6749 6653 6752
rect 6687 6780 6699 6783
rect 7190 6780 7196 6792
rect 6687 6752 7196 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 8312 6780 8340 6888
rect 8573 6851 8631 6857
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8619 6820 9045 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 9033 6817 9045 6820
rect 9079 6848 9091 6851
rect 9306 6848 9312 6860
rect 9079 6820 9312 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 10686 6808 10692 6860
rect 10744 6808 10750 6860
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11790 6848 11796 6860
rect 11296 6820 11796 6848
rect 11296 6808 11302 6820
rect 11790 6808 11796 6820
rect 11848 6848 11854 6860
rect 12345 6851 12403 6857
rect 12345 6848 12357 6851
rect 11848 6820 12357 6848
rect 11848 6808 11854 6820
rect 12345 6817 12357 6820
rect 12391 6817 12403 6851
rect 12345 6811 12403 6817
rect 12802 6808 12808 6860
rect 12860 6808 12866 6860
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8312 6752 8493 6780
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 10962 6780 10968 6792
rect 10827 6752 10968 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12526 6780 12532 6792
rect 12483 6752 12532 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12526 6740 12532 6752
rect 12584 6780 12590 6792
rect 13538 6780 13544 6792
rect 12584 6752 13544 6780
rect 12584 6740 12590 6752
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 6365 6715 6423 6721
rect 6365 6681 6377 6715
rect 6411 6681 6423 6715
rect 6365 6675 6423 6681
rect 6457 6715 6515 6721
rect 6457 6681 6469 6715
rect 6503 6712 6515 6715
rect 7466 6712 7472 6724
rect 6503 6684 7472 6712
rect 6503 6681 6515 6684
rect 6457 6675 6515 6681
rect 4356 6616 6224 6644
rect 6380 6644 6408 6675
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 7558 6644 7564 6656
rect 6380 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12894 6644 12900 6656
rect 12676 6616 12900 6644
rect 12676 6604 12682 6616
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 1104 6554 17756 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 17756 6554
rect 1104 6480 17756 6502
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3878 6440 3884 6452
rect 3191 6412 3884 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 7098 6440 7104 6452
rect 5920 6412 7104 6440
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 4890 6264 4896 6316
rect 4948 6264 4954 6316
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 5626 6264 5632 6316
rect 5684 6264 5690 6316
rect 5920 6313 5948 6412
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7466 6400 7472 6452
rect 7524 6400 7530 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 9122 6440 9128 6452
rect 7616 6412 9128 6440
rect 7616 6400 7622 6412
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 13814 6440 13820 6452
rect 11348 6412 13820 6440
rect 6270 6332 6276 6384
rect 6328 6372 6334 6384
rect 11238 6372 11244 6384
rect 6328 6344 7696 6372
rect 6328 6332 6334 6344
rect 6840 6313 6868 6344
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7558 6304 7564 6316
rect 6963 6276 7564 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 7668 6313 7696 6344
rect 11072 6344 11244 6372
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 8938 6304 8944 6316
rect 7699 6276 8944 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 11072 6313 11100 6344
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 11348 6381 11376 6412
rect 11333 6375 11391 6381
rect 11333 6341 11345 6375
rect 11379 6341 11391 6375
rect 11333 6335 11391 6341
rect 11790 6332 11796 6384
rect 11848 6332 11854 6384
rect 11992 6381 12020 6412
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 11977 6375 12035 6381
rect 11977 6341 11989 6375
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6372 13139 6375
rect 13541 6375 13599 6381
rect 13541 6372 13553 6375
rect 13127 6344 13553 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13541 6341 13553 6344
rect 13587 6341 13599 6375
rect 13541 6335 13599 6341
rect 14550 6332 14556 6384
rect 14608 6332 14614 6384
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 4663 6208 5181 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7190 6236 7196 6248
rect 7147 6208 7196 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 5813 6171 5871 6177
rect 5813 6137 5825 6171
rect 5859 6168 5871 6171
rect 7024 6168 7052 6199
rect 7190 6196 7196 6208
rect 7248 6236 7254 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7248 6208 7297 6236
rect 7248 6196 7254 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 9398 6236 9404 6248
rect 7524 6208 9404 6236
rect 7524 6196 7530 6208
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 7484 6168 7512 6196
rect 5859 6140 6960 6168
rect 7024 6140 7512 6168
rect 11164 6168 11192 6267
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 12802 6264 12808 6316
rect 12860 6264 12866 6316
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12345 6239 12403 6245
rect 12345 6236 12357 6239
rect 12308 6208 12357 6236
rect 12308 6196 12314 6208
rect 12345 6205 12357 6208
rect 12391 6205 12403 6239
rect 12345 6199 12403 6205
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 13078 6236 13084 6248
rect 12492 6208 13084 6236
rect 12492 6196 12498 6208
rect 13078 6196 13084 6208
rect 13136 6236 13142 6248
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 13136 6208 13277 6236
rect 13136 6196 13142 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 13596 6208 15301 6236
rect 13596 6196 13602 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 12526 6168 12532 6180
rect 11164 6140 12532 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 6638 6060 6644 6112
rect 6696 6060 6702 6112
rect 6932 6100 6960 6140
rect 7006 6100 7012 6112
rect 6932 6072 7012 6100
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7374 6060 7380 6112
rect 7432 6060 7438 6112
rect 11330 6060 11336 6112
rect 11388 6060 11394 6112
rect 11609 6103 11667 6109
rect 11609 6069 11621 6103
rect 11655 6100 11667 6103
rect 11698 6100 11704 6112
rect 11655 6072 11704 6100
rect 11655 6069 11667 6072
rect 11609 6063 11667 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11808 6109 11836 6140
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 11793 6103 11851 6109
rect 11793 6069 11805 6103
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 12437 6103 12495 6109
rect 12437 6069 12449 6103
rect 12483 6100 12495 6103
rect 12894 6100 12900 6112
rect 12483 6072 12900 6100
rect 12483 6069 12495 6072
rect 12437 6063 12495 6069
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 1104 6010 17756 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 17756 6010
rect 1104 5936 17756 5958
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 14550 5856 14556 5908
rect 14608 5856 14614 5908
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 11698 5828 11704 5840
rect 9180 5800 11704 5828
rect 9180 5788 9186 5800
rect 5721 5763 5779 5769
rect 5721 5729 5733 5763
rect 5767 5760 5779 5763
rect 6638 5760 6644 5772
rect 5767 5732 6644 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 9600 5769 9628 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5729 9643 5763
rect 9585 5723 9643 5729
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5760 9919 5763
rect 10318 5760 10324 5772
rect 9907 5732 10324 5760
rect 9907 5729 9919 5732
rect 9861 5723 9919 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 3844 5664 4077 5692
rect 3844 5652 3850 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 4080 5624 4108 5655
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 5905 5695 5963 5701
rect 5905 5692 5917 5695
rect 5868 5664 5917 5692
rect 5868 5652 5874 5664
rect 5905 5661 5917 5664
rect 5951 5692 5963 5695
rect 7374 5692 7380 5704
rect 5951 5664 7380 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11388 5664 11621 5692
rect 11388 5652 11394 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11698 5652 11704 5704
rect 11756 5692 11762 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11756 5664 11805 5692
rect 11756 5652 11762 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14645 5695 14703 5701
rect 14645 5692 14657 5695
rect 14332 5664 14657 5692
rect 14332 5652 14338 5664
rect 14645 5661 14657 5664
rect 14691 5692 14703 5695
rect 15102 5692 15108 5704
rect 14691 5664 15108 5692
rect 14691 5661 14703 5664
rect 14645 5655 14703 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 4080 5596 8432 5624
rect 8404 5568 8432 5596
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6638 5556 6644 5568
rect 6135 5528 6644 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 10962 5556 10968 5568
rect 8444 5528 10968 5556
rect 8444 5516 8450 5528
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 12342 5556 12348 5568
rect 11747 5528 12348 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 1104 5466 17756 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 17756 5466
rect 1104 5392 17756 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6822 5352 6828 5364
rect 5684 5324 6828 5352
rect 5684 5312 5690 5324
rect 6822 5312 6828 5324
rect 6880 5352 6886 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 6880 5324 8401 5352
rect 6880 5312 6886 5324
rect 8389 5321 8401 5324
rect 8435 5352 8447 5355
rect 10226 5352 10232 5364
rect 8435 5324 10232 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 10226 5312 10232 5324
rect 10284 5352 10290 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10284 5324 10517 5352
rect 10284 5312 10290 5324
rect 10505 5321 10517 5324
rect 10551 5352 10563 5355
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 10551 5324 12541 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 12529 5321 12541 5324
rect 12575 5352 12587 5355
rect 12618 5352 12624 5364
rect 12575 5324 12624 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 5592 5256 6776 5284
rect 5592 5244 5598 5256
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6748 5225 6776 5256
rect 7098 5244 7104 5296
rect 7156 5284 7162 5296
rect 7156 5256 10824 5284
rect 7156 5244 7162 5256
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5216 6791 5219
rect 6779 5188 6960 5216
rect 6779 5185 6791 5188
rect 6733 5179 6791 5185
rect 6932 5080 6960 5188
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8110 5216 8116 5228
rect 7064 5188 8116 5216
rect 7064 5176 7070 5188
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 8680 5225 8708 5256
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 7098 5108 7104 5160
rect 7156 5108 7162 5160
rect 8312 5148 8340 5179
rect 10318 5176 10324 5228
rect 10376 5176 10382 5228
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 10686 5216 10692 5228
rect 10459 5188 10692 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10428 5148 10456 5179
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 10796 5225 10824 5256
rect 10870 5244 10876 5296
rect 10928 5284 10934 5296
rect 12437 5287 12495 5293
rect 12437 5284 12449 5287
rect 10928 5256 12449 5284
rect 10928 5244 10934 5256
rect 12437 5253 12449 5256
rect 12483 5284 12495 5287
rect 12710 5284 12716 5296
rect 12483 5256 12716 5284
rect 12483 5253 12495 5256
rect 12437 5247 12495 5253
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 8312 5120 10456 5148
rect 10796 5148 10824 5179
rect 12342 5176 12348 5228
rect 12400 5176 12406 5228
rect 12250 5148 12256 5160
rect 10796 5120 12256 5148
rect 8312 5080 8340 5120
rect 12250 5108 12256 5120
rect 12308 5148 12314 5160
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 12308 5120 12817 5148
rect 12308 5108 12314 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 10689 5083 10747 5089
rect 10689 5080 10701 5083
rect 6932 5052 8340 5080
rect 8588 5052 10701 5080
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 6822 5012 6828 5024
rect 6411 4984 6828 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7926 4972 7932 5024
rect 7984 4972 7990 5024
rect 8110 4972 8116 5024
rect 8168 5012 8174 5024
rect 8588 5021 8616 5052
rect 10689 5049 10701 5052
rect 10735 5080 10747 5083
rect 12713 5083 12771 5089
rect 12713 5080 12725 5083
rect 10735 5052 12725 5080
rect 10735 5049 10747 5052
rect 10689 5043 10747 5049
rect 12713 5049 12725 5052
rect 12759 5080 12771 5083
rect 12894 5080 12900 5092
rect 12759 5052 12900 5080
rect 12759 5049 12771 5052
rect 12713 5043 12771 5049
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 8168 4984 8585 5012
rect 8168 4972 8174 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 8573 4975 8631 4981
rect 10045 5015 10103 5021
rect 10045 4981 10057 5015
rect 10091 5012 10103 5015
rect 10134 5012 10140 5024
rect 10091 4984 10140 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 12066 4972 12072 5024
rect 12124 4972 12130 5024
rect 1104 4922 17756 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 17756 4922
rect 1104 4848 17756 4870
rect 12066 4768 12072 4820
rect 12124 4808 12130 4820
rect 12326 4811 12384 4817
rect 12326 4808 12338 4811
rect 12124 4780 12338 4808
rect 12124 4768 12130 4780
rect 12326 4777 12338 4780
rect 12372 4777 12384 4811
rect 12326 4771 12384 4777
rect 13814 4768 13820 4820
rect 13872 4768 13878 4820
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 6546 4672 6552 4684
rect 5215 4644 6552 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 6972 4644 7205 4672
rect 6972 4632 6978 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 9861 4675 9919 4681
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 9907 4644 12081 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 12069 4641 12081 4644
rect 12115 4672 12127 4675
rect 13078 4672 13084 4684
rect 12115 4644 13084 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 8386 4564 8392 4616
rect 8444 4564 8450 4616
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 11480 4576 11897 4604
rect 11480 4564 11486 4576
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 11885 4567 11943 4573
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 6454 4496 6460 4548
rect 6512 4496 6518 4548
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 6917 4539 6975 4545
rect 6917 4536 6929 4539
rect 6880 4508 6929 4536
rect 6880 4496 6886 4508
rect 6917 4505 6929 4508
rect 6963 4505 6975 4539
rect 6917 4499 6975 4505
rect 10134 4496 10140 4548
rect 10192 4496 10198 4548
rect 11146 4496 11152 4548
rect 11204 4496 11210 4548
rect 14185 4539 14243 4545
rect 14185 4536 14197 4539
rect 13570 4508 14197 4536
rect 14185 4505 14197 4508
rect 14231 4505 14243 4539
rect 14185 4499 14243 4505
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8444 4440 8493 4468
rect 8444 4428 8450 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 1104 4378 17756 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 17756 4378
rect 1104 4304 17756 4326
rect 11057 4267 11115 4273
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11146 4264 11152 4276
rect 11103 4236 11152 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 7653 4199 7711 4205
rect 7653 4165 7665 4199
rect 7699 4196 7711 4199
rect 7926 4196 7932 4208
rect 7699 4168 7932 4196
rect 7699 4165 7711 4168
rect 7653 4159 7711 4165
rect 7926 4156 7932 4168
rect 7984 4156 7990 4208
rect 8386 4156 8392 4208
rect 8444 4156 8450 4208
rect 16574 4196 16580 4208
rect 14292 4168 16580 4196
rect 14292 4140 14320 4168
rect 16574 4156 16580 4168
rect 16632 4156 16638 4208
rect 6454 4088 6460 4140
rect 6512 4088 6518 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6564 4060 6592 4091
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 6972 4100 7389 4128
rect 6972 4088 6978 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 9398 4088 9404 4140
rect 9456 4088 9462 4140
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 11020 4100 11161 4128
rect 11020 4088 11026 4100
rect 11149 4097 11161 4100
rect 11195 4128 11207 4131
rect 14274 4128 14280 4140
rect 11195 4100 14280 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 8294 4060 8300 4072
rect 6564 4032 8300 4060
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 1104 3834 17756 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 17756 3834
rect 1104 3760 17756 3782
rect 16574 3544 16580 3596
rect 16632 3544 16638 3596
rect 17402 3476 17408 3528
rect 17460 3476 17466 3528
rect 1104 3290 17756 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 17756 3290
rect 1104 3216 17756 3238
rect 1104 2746 17756 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 17756 2746
rect 1104 2672 17756 2694
rect 1104 2202 17756 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 17756 2202
rect 1104 2128 17756 2150
<< via1 >>
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 7196 18411 7248 18420
rect 7196 18377 7205 18411
rect 7205 18377 7239 18411
rect 7239 18377 7248 18411
rect 7196 18368 7248 18377
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 11704 18411 11756 18420
rect 11704 18377 11713 18411
rect 11713 18377 11747 18411
rect 11747 18377 11756 18411
rect 11704 18368 11756 18377
rect 12992 18411 13044 18420
rect 12992 18377 13001 18411
rect 13001 18377 13035 18411
rect 13035 18377 13044 18411
rect 12992 18368 13044 18377
rect 10508 18343 10560 18352
rect 10508 18309 10517 18343
rect 10517 18309 10551 18343
rect 10551 18309 10560 18343
rect 10508 18300 10560 18309
rect 3884 18232 3936 18284
rect 6092 18275 6144 18284
rect 6092 18241 6101 18275
rect 6101 18241 6135 18275
rect 6135 18241 6144 18275
rect 6092 18232 6144 18241
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 7104 18232 7156 18284
rect 7748 18232 7800 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 10876 18232 10928 18284
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 13912 18164 13964 18216
rect 10692 18139 10744 18148
rect 10692 18105 10701 18139
rect 10701 18105 10735 18139
rect 10735 18105 10744 18139
rect 10692 18096 10744 18105
rect 2136 18028 2188 18080
rect 4528 18028 4580 18080
rect 6000 18028 6052 18080
rect 6920 18028 6972 18080
rect 9680 18028 9732 18080
rect 11520 18028 11572 18080
rect 12532 18071 12584 18080
rect 12532 18037 12541 18071
rect 12541 18037 12575 18071
rect 12575 18037 12584 18071
rect 12532 18028 12584 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 2350 17926 2402 17978
rect 2414 17926 2466 17978
rect 2478 17926 2530 17978
rect 2542 17926 2594 17978
rect 2606 17926 2658 17978
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 11888 17824 11940 17876
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 2780 17688 2832 17740
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 6368 17620 6420 17672
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 15660 17620 15712 17672
rect 2136 17552 2188 17604
rect 6000 17595 6052 17604
rect 2504 17484 2556 17536
rect 4068 17484 4120 17536
rect 6000 17561 6034 17595
rect 6034 17561 6052 17595
rect 6000 17552 6052 17561
rect 7840 17552 7892 17604
rect 9496 17595 9548 17604
rect 9496 17561 9530 17595
rect 9530 17561 9548 17595
rect 9496 17552 9548 17561
rect 10968 17595 11020 17604
rect 10968 17561 11002 17595
rect 11002 17561 11020 17595
rect 10968 17552 11020 17561
rect 11060 17552 11112 17604
rect 14924 17595 14976 17604
rect 14924 17561 14958 17595
rect 14958 17561 14976 17595
rect 4620 17484 4672 17536
rect 6460 17484 6512 17536
rect 8300 17484 8352 17536
rect 8668 17484 8720 17536
rect 10600 17527 10652 17536
rect 10600 17493 10609 17527
rect 10609 17493 10643 17527
rect 10643 17493 10652 17527
rect 14924 17552 14976 17561
rect 10600 17484 10652 17493
rect 16028 17527 16080 17536
rect 16028 17493 16037 17527
rect 16037 17493 16071 17527
rect 16071 17493 16080 17527
rect 16028 17484 16080 17493
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 1768 17280 1820 17332
rect 2504 17323 2556 17332
rect 2504 17289 2513 17323
rect 2513 17289 2547 17323
rect 2547 17289 2556 17323
rect 2504 17280 2556 17289
rect 4068 17280 4120 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 7840 17323 7892 17332
rect 7840 17289 7849 17323
rect 7849 17289 7883 17323
rect 7883 17289 7892 17323
rect 7840 17280 7892 17289
rect 10968 17280 11020 17332
rect 13912 17280 13964 17332
rect 5908 17212 5960 17264
rect 2228 17144 2280 17196
rect 3884 17187 3936 17196
rect 3884 17153 3893 17187
rect 3893 17153 3927 17187
rect 3927 17153 3936 17187
rect 3884 17144 3936 17153
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 6644 17187 6696 17196
rect 6644 17153 6678 17187
rect 6678 17153 6696 17187
rect 6644 17144 6696 17153
rect 6920 17144 6972 17196
rect 2136 17076 2188 17128
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 8300 17187 8352 17196
rect 8300 17153 8309 17187
rect 8309 17153 8343 17187
rect 8343 17153 8352 17187
rect 8300 17144 8352 17153
rect 9404 17144 9456 17196
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 9588 17144 9640 17196
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11888 17144 11940 17196
rect 14004 17144 14056 17196
rect 14280 17144 14332 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 16948 17076 17000 17128
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 13084 16940 13136 16992
rect 13820 17008 13872 17060
rect 15108 17008 15160 17060
rect 16764 17008 16816 17060
rect 14096 16940 14148 16992
rect 16580 16940 16632 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 2350 16838 2402 16890
rect 2414 16838 2466 16890
rect 2478 16838 2530 16890
rect 2542 16838 2594 16890
rect 2606 16838 2658 16890
rect 6644 16736 6696 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 8208 16736 8260 16788
rect 11888 16736 11940 16788
rect 4712 16668 4764 16720
rect 10968 16668 11020 16720
rect 7748 16600 7800 16652
rect 9496 16600 9548 16652
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16672 16600 16724 16652
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 9680 16532 9732 16584
rect 16580 16464 16632 16516
rect 14188 16396 14240 16448
rect 16948 16396 17000 16448
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 14924 16235 14976 16244
rect 14924 16201 14933 16235
rect 14933 16201 14967 16235
rect 14967 16201 14976 16235
rect 14924 16192 14976 16201
rect 14096 16167 14148 16176
rect 14096 16133 14105 16167
rect 14105 16133 14139 16167
rect 14139 16133 14148 16167
rect 14096 16124 14148 16133
rect 3884 16056 3936 16108
rect 5448 16056 5500 16108
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 14188 16099 14240 16108
rect 14188 16065 14197 16099
rect 14197 16065 14231 16099
rect 14231 16065 14240 16099
rect 14188 16056 14240 16065
rect 14556 16056 14608 16108
rect 15108 16099 15160 16108
rect 15108 16065 15117 16099
rect 15117 16065 15151 16099
rect 15151 16065 15160 16099
rect 15108 16056 15160 16065
rect 16028 16056 16080 16108
rect 14096 15988 14148 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 14464 15920 14516 15972
rect 2688 15895 2740 15904
rect 2688 15861 2697 15895
rect 2697 15861 2731 15895
rect 2731 15861 2740 15895
rect 2688 15852 2740 15861
rect 11336 15852 11388 15904
rect 12256 15852 12308 15904
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 2350 15750 2402 15802
rect 2414 15750 2466 15802
rect 2478 15750 2530 15802
rect 2542 15750 2594 15802
rect 2606 15750 2658 15802
rect 2872 15648 2924 15700
rect 6736 15648 6788 15700
rect 8024 15648 8076 15700
rect 10048 15648 10100 15700
rect 11980 15648 12032 15700
rect 7932 15580 7984 15632
rect 12532 15648 12584 15700
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 13912 15648 13964 15700
rect 14004 15580 14056 15632
rect 1400 15444 1452 15496
rect 2780 15512 2832 15564
rect 5908 15512 5960 15564
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 5448 15444 5500 15496
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6460 15487 6512 15496
rect 6460 15453 6467 15487
rect 6467 15453 6512 15487
rect 6460 15444 6512 15453
rect 6736 15487 6788 15496
rect 6736 15453 6769 15487
rect 6769 15453 6788 15487
rect 6736 15444 6788 15453
rect 6920 15444 6972 15496
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 7288 15512 7340 15564
rect 7564 15444 7616 15496
rect 7656 15444 7708 15496
rect 8116 15444 8168 15496
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 15660 15512 15712 15564
rect 11520 15444 11572 15453
rect 2688 15376 2740 15428
rect 4344 15376 4396 15428
rect 6184 15376 6236 15428
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 6828 15308 6880 15360
rect 7472 15308 7524 15360
rect 9036 15419 9088 15428
rect 9036 15385 9045 15419
rect 9045 15385 9079 15419
rect 9079 15385 9088 15419
rect 9036 15376 9088 15385
rect 9496 15376 9548 15428
rect 8024 15308 8076 15360
rect 9956 15308 10008 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 11980 15419 12032 15428
rect 11980 15385 11989 15419
rect 11989 15385 12023 15419
rect 12023 15385 12032 15419
rect 11980 15376 12032 15385
rect 12256 15376 12308 15428
rect 12624 15419 12676 15428
rect 12624 15385 12633 15419
rect 12633 15385 12667 15419
rect 12667 15385 12676 15419
rect 12624 15376 12676 15385
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 13636 15444 13688 15496
rect 13728 15376 13780 15428
rect 17224 15444 17276 15496
rect 15844 15376 15896 15428
rect 12900 15308 12952 15360
rect 13268 15308 13320 15360
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 1952 15104 2004 15156
rect 2872 15104 2924 15156
rect 4344 15104 4396 15156
rect 5540 15104 5592 15156
rect 6920 15147 6972 15156
rect 6920 15113 6929 15147
rect 6929 15113 6963 15147
rect 6963 15113 6972 15147
rect 6920 15104 6972 15113
rect 7012 15104 7064 15156
rect 9404 15104 9456 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 6736 15036 6788 15088
rect 7564 15036 7616 15088
rect 848 14968 900 15020
rect 2228 14968 2280 15020
rect 4528 14968 4580 15020
rect 6920 14968 6972 15020
rect 7748 14968 7800 15020
rect 2320 14900 2372 14952
rect 4436 14832 4488 14884
rect 6000 14900 6052 14952
rect 6276 14900 6328 14952
rect 7012 14900 7064 14952
rect 7104 14900 7156 14952
rect 7656 14900 7708 14952
rect 8116 15036 8168 15088
rect 11336 15104 11388 15156
rect 11428 15104 11480 15156
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 9956 14968 10008 15020
rect 13084 15104 13136 15156
rect 14740 15104 14792 15156
rect 15844 15147 15896 15156
rect 15844 15113 15853 15147
rect 15853 15113 15887 15147
rect 15887 15113 15896 15147
rect 15844 15104 15896 15113
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 13268 15036 13320 15088
rect 13084 14968 13136 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 5448 14764 5500 14816
rect 9956 14764 10008 14816
rect 11152 14832 11204 14884
rect 13544 14900 13596 14952
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 15200 14900 15252 14952
rect 16120 14900 16172 14952
rect 17316 14900 17368 14952
rect 14924 14832 14976 14884
rect 12808 14764 12860 14816
rect 2350 14662 2402 14714
rect 2414 14662 2466 14714
rect 2478 14662 2530 14714
rect 2542 14662 2594 14714
rect 2606 14662 2658 14714
rect 6552 14560 6604 14612
rect 12900 14560 12952 14612
rect 17040 14560 17092 14612
rect 6460 14492 6512 14544
rect 7564 14492 7616 14544
rect 6184 14424 6236 14476
rect 5448 14356 5500 14408
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 6092 14399 6144 14408
rect 6092 14365 6102 14399
rect 6102 14365 6136 14399
rect 6136 14365 6144 14399
rect 7472 14424 7524 14476
rect 12624 14424 12676 14476
rect 14556 14424 14608 14476
rect 6092 14356 6144 14365
rect 6736 14356 6788 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 6368 14331 6420 14340
rect 6368 14297 6377 14331
rect 6377 14297 6411 14331
rect 6411 14297 6420 14331
rect 6368 14288 6420 14297
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 4252 14220 4304 14272
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 1400 14016 1452 14068
rect 2412 13948 2464 14000
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 8392 14016 8444 14068
rect 9312 14016 9364 14068
rect 11704 14016 11756 14068
rect 12900 14016 12952 14068
rect 14372 14059 14424 14068
rect 14372 14025 14381 14059
rect 14381 14025 14415 14059
rect 14415 14025 14424 14059
rect 14372 14016 14424 14025
rect 4252 13948 4304 14000
rect 9404 13948 9456 14000
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 4528 13880 4580 13932
rect 5448 13880 5500 13932
rect 7932 13923 7984 13932
rect 7932 13889 7966 13923
rect 7966 13889 7984 13923
rect 7932 13880 7984 13889
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 11336 13948 11388 14000
rect 10784 13923 10836 13932
rect 10784 13889 10791 13923
rect 10791 13889 10836 13923
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 3516 13812 3568 13864
rect 3700 13855 3752 13864
rect 3700 13821 3709 13855
rect 3709 13821 3743 13855
rect 3743 13821 3752 13855
rect 3700 13812 3752 13821
rect 6184 13812 6236 13864
rect 6552 13744 6604 13796
rect 7104 13812 7156 13864
rect 7656 13855 7708 13864
rect 7656 13821 7665 13855
rect 7665 13821 7699 13855
rect 7699 13821 7708 13855
rect 7656 13812 7708 13821
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10048 13812 10100 13821
rect 10784 13880 10836 13889
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11152 13880 11204 13932
rect 13268 13880 13320 13932
rect 14280 13880 14332 13932
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 14648 13923 14700 13932
rect 14648 13889 14655 13923
rect 14655 13889 14700 13923
rect 14648 13880 14700 13889
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 11796 13676 11848 13728
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 14924 13923 14976 13932
rect 14924 13889 14938 13923
rect 14938 13889 14972 13923
rect 14972 13889 14976 13923
rect 17224 14059 17276 14068
rect 17224 14025 17233 14059
rect 17233 14025 17267 14059
rect 17267 14025 17276 14059
rect 17224 14016 17276 14025
rect 14924 13880 14976 13889
rect 16120 13923 16172 13932
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 13820 13744 13872 13796
rect 17224 13812 17276 13864
rect 14004 13744 14056 13796
rect 14556 13744 14608 13796
rect 16304 13744 16356 13796
rect 15752 13719 15804 13728
rect 15752 13685 15761 13719
rect 15761 13685 15795 13719
rect 15795 13685 15804 13719
rect 15752 13676 15804 13685
rect 2350 13574 2402 13626
rect 2414 13574 2466 13626
rect 2478 13574 2530 13626
rect 2542 13574 2594 13626
rect 2606 13574 2658 13626
rect 1676 13472 1728 13524
rect 3700 13472 3752 13524
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 13268 13515 13320 13524
rect 13268 13481 13277 13515
rect 13277 13481 13311 13515
rect 13311 13481 13320 13515
rect 13268 13472 13320 13481
rect 16028 13472 16080 13524
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 2136 13336 2188 13388
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 8392 13379 8444 13388
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 13268 13336 13320 13388
rect 15660 13336 15712 13388
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 848 13268 900 13320
rect 3332 13268 3384 13320
rect 5724 13268 5776 13320
rect 7012 13268 7064 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 14464 13311 14516 13320
rect 14464 13277 14471 13311
rect 14471 13277 14516 13311
rect 14464 13268 14516 13277
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 14924 13268 14976 13320
rect 15752 13268 15804 13320
rect 4528 13200 4580 13252
rect 7380 13243 7432 13252
rect 7380 13209 7389 13243
rect 7389 13209 7423 13243
rect 7423 13209 7432 13243
rect 7380 13200 7432 13209
rect 9312 13243 9364 13252
rect 9312 13209 9321 13243
rect 9321 13209 9355 13243
rect 9355 13209 9364 13243
rect 9312 13200 9364 13209
rect 10048 13200 10100 13252
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 12532 13200 12584 13252
rect 14648 13243 14700 13252
rect 14648 13209 14657 13243
rect 14657 13209 14691 13243
rect 14691 13209 14700 13243
rect 14648 13200 14700 13209
rect 3516 13132 3568 13184
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 3516 12928 3568 12980
rect 6092 12928 6144 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 9312 12928 9364 12980
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 5724 12903 5776 12912
rect 5724 12869 5733 12903
rect 5733 12869 5767 12903
rect 5767 12869 5776 12903
rect 5724 12860 5776 12869
rect 6276 12860 6328 12912
rect 7104 12860 7156 12912
rect 6000 12792 6052 12844
rect 6460 12835 6512 12844
rect 6460 12801 6470 12835
rect 6470 12801 6504 12835
rect 6504 12801 6512 12835
rect 6460 12792 6512 12801
rect 6828 12835 6880 12844
rect 6828 12801 6861 12835
rect 6861 12801 6880 12835
rect 6828 12792 6880 12801
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10784 12792 10836 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 13360 12792 13412 12844
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 14188 12792 14240 12844
rect 15016 12792 15068 12844
rect 17224 12860 17276 12912
rect 17408 12835 17460 12844
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 5540 12724 5592 12776
rect 5724 12724 5776 12776
rect 10876 12724 10928 12776
rect 14924 12724 14976 12776
rect 4252 12656 4304 12708
rect 6460 12656 6512 12708
rect 13636 12699 13688 12708
rect 13636 12665 13645 12699
rect 13645 12665 13679 12699
rect 13679 12665 13688 12699
rect 13636 12656 13688 12665
rect 13820 12656 13872 12708
rect 4528 12588 4580 12640
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 2350 12486 2402 12538
rect 2414 12486 2466 12538
rect 2478 12486 2530 12538
rect 2542 12486 2594 12538
rect 2606 12486 2658 12538
rect 2872 12384 2924 12436
rect 4252 12384 4304 12436
rect 5632 12384 5684 12436
rect 6184 12384 6236 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 5356 12316 5408 12368
rect 5540 12316 5592 12368
rect 5816 12316 5868 12368
rect 5908 12316 5960 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 4344 12180 4396 12232
rect 7840 12316 7892 12368
rect 7932 12359 7984 12368
rect 7932 12325 7941 12359
rect 7941 12325 7975 12359
rect 7975 12325 7984 12359
rect 7932 12316 7984 12325
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 4896 12180 4948 12232
rect 5264 12180 5316 12232
rect 5540 12223 5592 12232
rect 5540 12189 5548 12223
rect 5548 12189 5582 12223
rect 5582 12189 5592 12223
rect 5540 12180 5592 12189
rect 6000 12223 6052 12232
rect 6000 12189 6008 12223
rect 6008 12189 6042 12223
rect 6042 12189 6052 12223
rect 6000 12180 6052 12189
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 7196 12180 7248 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 8208 12223 8260 12232
rect 8208 12189 8217 12223
rect 8217 12189 8251 12223
rect 8251 12189 8260 12223
rect 8208 12180 8260 12189
rect 4252 12044 4304 12096
rect 4620 12044 4672 12096
rect 5080 12044 5132 12096
rect 5632 12044 5684 12096
rect 6184 12112 6236 12164
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 7472 12044 7524 12096
rect 7840 12044 7892 12096
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 10784 12180 10836 12232
rect 15016 12384 15068 12436
rect 14464 12248 14516 12300
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 15844 12180 15896 12232
rect 14556 12112 14608 12164
rect 16764 12248 16816 12300
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 16856 12180 16908 12189
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 14740 12044 14792 12096
rect 15936 12044 15988 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 1676 11840 1728 11892
rect 2872 11840 2924 11892
rect 5264 11883 5316 11892
rect 5264 11849 5273 11883
rect 5273 11849 5307 11883
rect 5307 11849 5316 11883
rect 5264 11840 5316 11849
rect 5356 11840 5408 11892
rect 6184 11840 6236 11892
rect 7288 11840 7340 11892
rect 7932 11840 7984 11892
rect 15568 11840 15620 11892
rect 2688 11772 2740 11824
rect 2136 11704 2188 11756
rect 4344 11704 4396 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 5540 11772 5592 11824
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 4620 11636 4672 11688
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 5816 11747 5868 11756
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6460 11704 6512 11756
rect 14740 11772 14792 11824
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 10600 11704 10652 11756
rect 11428 11636 11480 11688
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 16120 11704 16172 11756
rect 17316 11704 17368 11756
rect 12900 11636 12952 11688
rect 14188 11636 14240 11688
rect 14924 11636 14976 11688
rect 16764 11636 16816 11688
rect 17408 11611 17460 11620
rect 17408 11577 17417 11611
rect 17417 11577 17451 11611
rect 17451 11577 17460 11611
rect 17408 11568 17460 11577
rect 4068 11543 4120 11552
rect 4068 11509 4077 11543
rect 4077 11509 4111 11543
rect 4111 11509 4120 11543
rect 4068 11500 4120 11509
rect 4528 11500 4580 11552
rect 11980 11543 12032 11552
rect 11980 11509 11989 11543
rect 11989 11509 12023 11543
rect 12023 11509 12032 11543
rect 11980 11500 12032 11509
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 2350 11398 2402 11450
rect 2414 11398 2466 11450
rect 2478 11398 2530 11450
rect 2542 11398 2594 11450
rect 2606 11398 2658 11450
rect 5816 11296 5868 11348
rect 6092 11296 6144 11348
rect 7748 11296 7800 11348
rect 12624 11296 12676 11348
rect 12808 11339 12860 11348
rect 12808 11305 12817 11339
rect 12817 11305 12851 11339
rect 12851 11305 12860 11339
rect 12808 11296 12860 11305
rect 16488 11296 16540 11348
rect 11060 11160 11112 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 11980 11092 12032 11144
rect 15936 11203 15988 11212
rect 15936 11169 15945 11203
rect 15945 11169 15979 11203
rect 15979 11169 15988 11203
rect 15936 11160 15988 11169
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 10692 11024 10744 11076
rect 12072 11024 12124 11076
rect 12716 11092 12768 11144
rect 12808 11092 12860 11144
rect 13728 11092 13780 11144
rect 15568 11092 15620 11144
rect 2688 10956 2740 11008
rect 4528 10956 4580 11008
rect 9036 10956 9088 11008
rect 14464 11024 14516 11076
rect 16948 11024 17000 11076
rect 12440 10956 12492 11008
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 2688 10752 2740 10804
rect 5264 10752 5316 10804
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 7380 10752 7432 10804
rect 11796 10752 11848 10804
rect 13636 10752 13688 10804
rect 14832 10752 14884 10804
rect 16120 10795 16172 10804
rect 16120 10761 16129 10795
rect 16129 10761 16163 10795
rect 16163 10761 16172 10795
rect 16120 10752 16172 10761
rect 1308 10684 1360 10736
rect 10692 10727 10744 10736
rect 10692 10693 10701 10727
rect 10701 10693 10735 10727
rect 10735 10693 10744 10727
rect 10692 10684 10744 10693
rect 3148 10616 3200 10668
rect 2228 10548 2280 10600
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 4436 10616 4488 10668
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 5356 10659 5408 10668
rect 5356 10625 5395 10659
rect 5395 10625 5408 10659
rect 5356 10616 5408 10625
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 5908 10616 5960 10668
rect 6920 10616 6972 10668
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 5540 10480 5592 10532
rect 6000 10480 6052 10532
rect 1676 10412 1728 10464
rect 3516 10412 3568 10464
rect 3976 10412 4028 10464
rect 5356 10412 5408 10464
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 9956 10616 10008 10668
rect 10876 10616 10928 10668
rect 11244 10616 11296 10668
rect 7196 10480 7248 10532
rect 7748 10480 7800 10532
rect 8116 10480 8168 10532
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 8300 10412 8352 10464
rect 11980 10412 12032 10464
rect 12900 10412 12952 10464
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 14004 10412 14056 10464
rect 15108 10412 15160 10464
rect 15844 10412 15896 10464
rect 2350 10310 2402 10362
rect 2414 10310 2466 10362
rect 2478 10310 2530 10362
rect 2542 10310 2594 10362
rect 2606 10310 2658 10362
rect 5540 10208 5592 10260
rect 7472 10208 7524 10260
rect 7748 10208 7800 10260
rect 10968 10251 11020 10260
rect 10968 10217 10977 10251
rect 10977 10217 11011 10251
rect 11011 10217 11020 10251
rect 10968 10208 11020 10217
rect 16212 10208 16264 10260
rect 3792 10183 3844 10192
rect 3792 10149 3801 10183
rect 3801 10149 3835 10183
rect 3835 10149 3844 10183
rect 3792 10140 3844 10149
rect 2872 10072 2924 10124
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4528 10004 4580 10056
rect 5080 10004 5132 10056
rect 5908 10072 5960 10124
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 5724 10004 5776 10056
rect 7288 10072 7340 10124
rect 7564 10072 7616 10124
rect 6920 10004 6972 10056
rect 8024 10004 8076 10056
rect 10968 10072 11020 10124
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 13820 10072 13872 10124
rect 15016 10072 15068 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 15568 10047 15620 10056
rect 15568 10013 15577 10047
rect 15577 10013 15611 10047
rect 15611 10013 15620 10047
rect 15568 10004 15620 10013
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 9128 9936 9180 9988
rect 16580 9936 16632 9988
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3884 9868 3936 9920
rect 4436 9868 4488 9920
rect 5632 9868 5684 9920
rect 11336 9911 11388 9920
rect 11336 9877 11345 9911
rect 11345 9877 11379 9911
rect 11379 9877 11388 9911
rect 11336 9868 11388 9877
rect 11796 9868 11848 9920
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 3884 9664 3936 9716
rect 5908 9664 5960 9716
rect 6920 9664 6972 9716
rect 7656 9664 7708 9716
rect 7380 9596 7432 9648
rect 9312 9596 9364 9648
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10968 9528 11020 9580
rect 11060 9528 11112 9580
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 12440 9596 12492 9648
rect 16580 9596 16632 9648
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 9588 9435 9640 9444
rect 9588 9401 9597 9435
rect 9597 9401 9631 9435
rect 9631 9401 9640 9435
rect 9588 9392 9640 9401
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 11428 9460 11480 9512
rect 13912 9460 13964 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 16764 9460 16816 9512
rect 11336 9392 11388 9444
rect 13544 9392 13596 9444
rect 14648 9392 14700 9444
rect 16396 9392 16448 9444
rect 12532 9324 12584 9376
rect 12716 9324 12768 9376
rect 2350 9222 2402 9274
rect 2414 9222 2466 9274
rect 2478 9222 2530 9274
rect 2542 9222 2594 9274
rect 2606 9222 2658 9274
rect 9220 9120 9272 9172
rect 9312 9120 9364 9172
rect 10232 9120 10284 9172
rect 12992 9120 13044 9172
rect 3976 9052 4028 9104
rect 9864 9052 9916 9104
rect 12716 9095 12768 9104
rect 12716 9061 12725 9095
rect 12725 9061 12759 9095
rect 12759 9061 12768 9095
rect 12716 9052 12768 9061
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 3884 8916 3936 8925
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 6644 8984 6696 9036
rect 3884 8780 3936 8832
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 7472 8984 7524 9036
rect 7748 8984 7800 9036
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 4804 8848 4856 8900
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 7196 8916 7248 8968
rect 8116 8916 8168 8968
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 10784 8984 10836 9036
rect 12440 8984 12492 9036
rect 8300 8916 8352 8925
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 14004 9052 14056 9104
rect 4528 8780 4580 8832
rect 8024 8848 8076 8900
rect 10140 8848 10192 8900
rect 7012 8780 7064 8832
rect 12808 8780 12860 8832
rect 16304 8984 16356 9036
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 16396 8959 16448 8968
rect 16396 8925 16405 8959
rect 16405 8925 16439 8959
rect 16439 8925 16448 8959
rect 16396 8916 16448 8925
rect 13544 8848 13596 8900
rect 14556 8780 14608 8832
rect 15844 8780 15896 8832
rect 15936 8780 15988 8832
rect 16764 8780 16816 8832
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 2872 8508 2924 8560
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 3516 8372 3568 8424
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4528 8483 4580 8492
rect 4528 8449 4537 8483
rect 4537 8449 4571 8483
rect 4571 8449 4580 8483
rect 4528 8440 4580 8449
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5724 8576 5776 8628
rect 5448 8440 5500 8492
rect 5908 8440 5960 8492
rect 7932 8576 7984 8628
rect 12624 8576 12676 8628
rect 5540 8372 5592 8424
rect 5724 8372 5776 8424
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 7012 8440 7064 8492
rect 11428 8508 11480 8560
rect 7840 8440 7892 8492
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 11336 8440 11388 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13912 8483 13964 8492
rect 8208 8372 8260 8424
rect 5816 8304 5868 8356
rect 6552 8304 6604 8356
rect 6828 8304 6880 8356
rect 12624 8347 12676 8356
rect 12624 8313 12633 8347
rect 12633 8313 12667 8347
rect 12667 8313 12676 8347
rect 12624 8304 12676 8313
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 13912 8449 13920 8483
rect 13920 8449 13954 8483
rect 13954 8449 13964 8483
rect 13912 8440 13964 8449
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 16764 8372 16816 8424
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 1584 8236 1636 8288
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 8024 8236 8076 8288
rect 2350 8134 2402 8186
rect 2414 8134 2466 8186
rect 2478 8134 2530 8186
rect 2542 8134 2594 8186
rect 2606 8134 2658 8186
rect 1308 8032 1360 8084
rect 13176 8032 13228 8084
rect 16764 8032 16816 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 12624 7964 12676 8016
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 11336 7896 11388 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 3884 7871 3936 7880
rect 3884 7837 3893 7871
rect 3893 7837 3927 7871
rect 3927 7837 3936 7871
rect 3884 7828 3936 7837
rect 3976 7871 4028 7880
rect 3976 7837 3986 7871
rect 3986 7837 4020 7871
rect 4020 7837 4028 7871
rect 3976 7828 4028 7837
rect 7012 7828 7064 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 10232 7828 10284 7880
rect 11428 7828 11480 7880
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 11980 7760 12032 7812
rect 16764 7760 16816 7812
rect 848 7692 900 7744
rect 9588 7692 9640 7744
rect 10784 7692 10836 7744
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 1860 7488 1912 7540
rect 8116 7488 8168 7540
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 2228 7420 2280 7472
rect 2872 7420 2924 7472
rect 11060 7488 11112 7540
rect 12440 7488 12492 7540
rect 4896 7352 4948 7404
rect 7472 7352 7524 7404
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 11244 7420 11296 7472
rect 3792 7284 3844 7336
rect 10692 7352 10744 7404
rect 15568 7488 15620 7540
rect 15844 7488 15896 7540
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 14556 7463 14608 7472
rect 14556 7429 14565 7463
rect 14565 7429 14599 7463
rect 14599 7429 14608 7463
rect 14556 7420 14608 7429
rect 16856 7395 16908 7404
rect 9588 7284 9640 7336
rect 11428 7284 11480 7336
rect 15200 7284 15252 7336
rect 16856 7361 16865 7395
rect 16865 7361 16899 7395
rect 16899 7361 16908 7395
rect 16856 7352 16908 7361
rect 8944 7148 8996 7200
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 8208 6944 8260 6996
rect 2228 6808 2280 6860
rect 5632 6876 5684 6928
rect 3424 6740 3476 6792
rect 3792 6740 3844 6792
rect 3884 6740 3936 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 8208 6808 8260 6860
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 6552 6740 6604 6792
rect 7196 6740 7248 6792
rect 9312 6808 9364 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 11244 6808 11296 6860
rect 11796 6808 11848 6860
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 10968 6740 11020 6792
rect 12532 6740 12584 6792
rect 13544 6740 13596 6792
rect 7472 6672 7524 6724
rect 7564 6604 7616 6656
rect 12624 6604 12676 6656
rect 12900 6604 12952 6656
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 3884 6400 3936 6452
rect 3976 6332 4028 6384
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 7104 6400 7156 6452
rect 7472 6443 7524 6452
rect 7472 6409 7481 6443
rect 7481 6409 7515 6443
rect 7515 6409 7524 6443
rect 7472 6400 7524 6409
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 9128 6400 9180 6452
rect 6276 6332 6328 6384
rect 7564 6264 7616 6316
rect 8944 6264 8996 6316
rect 11244 6332 11296 6384
rect 11796 6375 11848 6384
rect 11796 6341 11805 6375
rect 11805 6341 11839 6375
rect 11839 6341 11848 6375
rect 11796 6332 11848 6341
rect 13820 6400 13872 6452
rect 14556 6332 14608 6384
rect 7196 6196 7248 6248
rect 7472 6196 7524 6248
rect 9404 6196 9456 6248
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 12256 6196 12308 6248
rect 12440 6196 12492 6248
rect 13084 6196 13136 6248
rect 13544 6196 13596 6248
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 7012 6060 7064 6112
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 11704 6060 11756 6112
rect 12532 6128 12584 6180
rect 12900 6060 12952 6112
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 9128 5788 9180 5840
rect 6644 5720 6696 5772
rect 11704 5788 11756 5840
rect 10324 5720 10376 5772
rect 3792 5652 3844 5704
rect 5816 5652 5868 5704
rect 7380 5652 7432 5704
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 11336 5652 11388 5704
rect 11704 5652 11756 5704
rect 14280 5652 14332 5704
rect 15108 5652 15160 5704
rect 6644 5516 6696 5568
rect 8392 5516 8444 5568
rect 10968 5516 11020 5568
rect 12348 5516 12400 5568
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 5632 5312 5684 5364
rect 6828 5355 6880 5364
rect 6828 5321 6837 5355
rect 6837 5321 6871 5355
rect 6871 5321 6880 5355
rect 6828 5312 6880 5321
rect 10232 5312 10284 5364
rect 12624 5312 12676 5364
rect 5540 5244 5592 5296
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7104 5244 7156 5296
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 8116 5176 8168 5228
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 10692 5176 10744 5228
rect 10876 5244 10928 5296
rect 12716 5244 12768 5296
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 12256 5108 12308 5160
rect 6828 4972 6880 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8116 4972 8168 5024
rect 12900 5040 12952 5092
rect 10140 4972 10192 5024
rect 12072 5015 12124 5024
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 12072 4768 12124 4820
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 6552 4632 6604 4684
rect 6920 4632 6972 4684
rect 13084 4632 13136 4684
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 11428 4564 11480 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 6460 4496 6512 4548
rect 6828 4496 6880 4548
rect 10140 4539 10192 4548
rect 10140 4505 10149 4539
rect 10149 4505 10183 4539
rect 10183 4505 10192 4539
rect 10140 4496 10192 4505
rect 11152 4496 11204 4548
rect 8392 4428 8444 4480
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 11152 4224 11204 4276
rect 7932 4156 7984 4208
rect 8392 4156 8444 4208
rect 16580 4156 16632 4208
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6920 4088 6972 4140
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 10968 4088 11020 4140
rect 14280 4088 14332 4140
rect 8300 4020 8352 4072
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
<< metal2 >>
rect 5814 20346 5870 21033
rect 7102 20346 7158 21033
rect 7746 20346 7802 21033
rect 8390 20346 8446 21033
rect 9034 20346 9090 21033
rect 9678 20346 9734 21033
rect 10322 20346 10378 21033
rect 10966 20346 11022 21033
rect 5814 20318 6132 20346
rect 5814 20233 5870 20318
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 6104 18290 6132 20318
rect 7102 20318 7236 20346
rect 7102 20233 7158 20318
rect 7208 18426 7236 20318
rect 7746 20318 7880 20346
rect 7746 20233 7802 20318
rect 7852 18426 7880 20318
rect 8390 20318 8524 20346
rect 8390 20233 8446 20318
rect 8496 18426 8524 20318
rect 9034 20318 9168 20346
rect 9034 20233 9090 20318
rect 9140 18426 9168 20318
rect 9678 20318 9996 20346
rect 9678 20233 9734 20318
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9968 18290 9996 20318
rect 10322 20318 10548 20346
rect 10322 20233 10378 20318
rect 10520 18358 10548 20318
rect 10888 20318 11022 20346
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10888 18290 10916 20318
rect 10966 20233 11022 20318
rect 11610 20346 11666 21033
rect 12254 20346 12310 21033
rect 12898 20346 12954 21033
rect 13542 20346 13598 21033
rect 11610 20318 11744 20346
rect 11610 20233 11666 20318
rect 11716 18426 11744 20318
rect 12254 20318 12388 20346
rect 12254 20233 12310 20318
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 12360 18290 12388 20318
rect 12898 20318 13032 20346
rect 12898 20233 12954 20318
rect 13004 18426 13032 20318
rect 13542 20318 13676 20346
rect 13542 20233 13598 20318
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13648 18290 13676 20318
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17338 1808 17614
rect 2148 17610 2176 18022
rect 2350 17980 2658 17989
rect 2350 17978 2356 17980
rect 2412 17978 2436 17980
rect 2492 17978 2516 17980
rect 2572 17978 2596 17980
rect 2652 17978 2658 17980
rect 2412 17926 2414 17978
rect 2594 17926 2596 17978
rect 2350 17924 2356 17926
rect 2412 17924 2436 17926
rect 2492 17924 2516 17926
rect 2572 17924 2596 17926
rect 2652 17924 2658 17926
rect 2350 17915 2658 17924
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2516 17338 2544 17478
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 17128 2188 17134
rect 1306 17096 1362 17105
rect 2136 17070 2188 17076
rect 1306 17031 1362 17040
rect 848 15020 900 15026
rect 848 14962 900 14968
rect 860 14929 888 14962
rect 846 14920 902 14929
rect 846 14855 902 14864
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 1320 10742 1348 17031
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1412 14074 1440 15438
rect 1964 15162 1992 15438
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 1412 13870 1440 14010
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1412 12306 1440 13806
rect 1688 13530 1716 13806
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 2148 13394 2176 17070
rect 2240 15026 2268 17138
rect 2350 16892 2658 16901
rect 2350 16890 2356 16892
rect 2412 16890 2436 16892
rect 2492 16890 2516 16892
rect 2572 16890 2596 16892
rect 2652 16890 2658 16892
rect 2412 16838 2414 16890
rect 2594 16838 2596 16890
rect 2350 16836 2356 16838
rect 2412 16836 2436 16838
rect 2492 16836 2516 16838
rect 2572 16836 2596 16838
rect 2652 16836 2658 16838
rect 2350 16827 2658 16836
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2350 15804 2658 15813
rect 2350 15802 2356 15804
rect 2412 15802 2436 15804
rect 2492 15802 2516 15804
rect 2572 15802 2596 15804
rect 2652 15802 2658 15804
rect 2412 15750 2414 15802
rect 2594 15750 2596 15802
rect 2350 15748 2356 15750
rect 2412 15748 2436 15750
rect 2492 15748 2516 15750
rect 2572 15748 2596 15750
rect 2652 15748 2658 15750
rect 2350 15739 2658 15748
rect 2700 15434 2728 15846
rect 2792 15570 2820 17682
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 3896 17202 3924 18226
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17338 4108 17478
rect 4172 17338 4200 17614
rect 4540 17338 4568 18022
rect 6012 17610 6040 18022
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6000 17604 6052 17610
rect 6000 17546 6052 17552
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4632 17338 4660 17478
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 3896 16114 3924 17138
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2884 15162 2912 15642
rect 4344 15428 4396 15434
rect 4344 15370 4396 15376
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 4356 15162 4384 15370
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4540 15026 4568 17274
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16726 4752 17070
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15502 5488 16050
rect 5920 15570 5948 17206
rect 6380 17202 6408 17614
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 2320 14952 2372 14958
rect 2240 14900 2320 14906
rect 2240 14894 2372 14900
rect 2240 14878 2360 14894
rect 4436 14884 4488 14890
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11898 1716 12106
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 2148 11762 2176 13330
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1308 10736 1360 10742
rect 1308 10678 1360 10684
rect 2240 10606 2268 14878
rect 4436 14826 4488 14832
rect 2350 14716 2658 14725
rect 2350 14714 2356 14716
rect 2412 14714 2436 14716
rect 2492 14714 2516 14716
rect 2572 14714 2596 14716
rect 2652 14714 2658 14716
rect 2412 14662 2414 14714
rect 2594 14662 2596 14714
rect 2350 14660 2356 14662
rect 2412 14660 2436 14662
rect 2492 14660 2516 14662
rect 2572 14660 2596 14662
rect 2652 14660 2658 14662
rect 2350 14651 2658 14660
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 2424 14006 2452 14214
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 4264 14006 4292 14214
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 2350 13628 2658 13637
rect 2350 13626 2356 13628
rect 2412 13626 2436 13628
rect 2492 13626 2516 13628
rect 2572 13626 2596 13628
rect 2652 13626 2658 13628
rect 2412 13574 2414 13626
rect 2594 13574 2596 13626
rect 2350 13572 2356 13574
rect 2412 13572 2436 13574
rect 2492 13572 2516 13574
rect 2572 13572 2596 13574
rect 2652 13572 2658 13574
rect 2350 13563 2658 13572
rect 3344 13326 3372 13874
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3528 13190 3556 13806
rect 3712 13530 3740 13806
rect 3700 13524 3752 13530
rect 3700 13466 3752 13472
rect 4448 13394 4476 14826
rect 5460 14822 5488 15438
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 15162 5580 15302
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 14414 5488 14758
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4540 13258 4568 13874
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 3528 12986 3556 13126
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 2350 12540 2658 12549
rect 2350 12538 2356 12540
rect 2412 12538 2436 12540
rect 2492 12538 2516 12540
rect 2572 12538 2596 12540
rect 2652 12538 2658 12540
rect 2412 12486 2414 12538
rect 2594 12486 2596 12538
rect 2350 12484 2356 12486
rect 2412 12484 2436 12486
rect 2492 12484 2516 12486
rect 2572 12484 2596 12486
rect 2652 12484 2658 12486
rect 2350 12475 2658 12484
rect 4264 12442 4292 12650
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 2884 11898 2912 12378
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2350 11452 2658 11461
rect 2350 11450 2356 11452
rect 2412 11450 2436 11452
rect 2492 11450 2516 11452
rect 2572 11450 2596 11452
rect 2652 11450 2658 11452
rect 2412 11398 2414 11450
rect 2594 11398 2596 11450
rect 2350 11396 2356 11398
rect 2412 11396 2436 11398
rect 2492 11396 2516 11398
rect 2572 11396 2596 11398
rect 2652 11396 2658 11398
rect 2350 11387 2658 11396
rect 2700 11014 2728 11766
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2700 10810 2728 10950
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 9994 1716 10406
rect 2350 10364 2658 10373
rect 2350 10362 2356 10364
rect 2412 10362 2436 10364
rect 2492 10362 2516 10364
rect 2572 10362 2596 10364
rect 2652 10362 2658 10364
rect 2412 10310 2414 10362
rect 2594 10310 2596 10362
rect 2350 10308 2356 10310
rect 2412 10308 2436 10310
rect 2492 10308 2516 10310
rect 2572 10308 2596 10310
rect 2652 10308 2658 10310
rect 2350 10299 2658 10308
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 1676 9988 1728 9994
rect 1676 9930 1728 9936
rect 2350 9276 2658 9285
rect 2350 9274 2356 9276
rect 2412 9274 2436 9276
rect 2492 9274 2516 9276
rect 2572 9274 2596 9276
rect 2652 9274 2658 9276
rect 2412 9222 2414 9274
rect 2594 9222 2596 9274
rect 2350 9220 2356 9222
rect 2412 9220 2436 9222
rect 2492 9220 2516 9222
rect 2572 9220 2596 9222
rect 2652 9220 2658 9222
rect 2350 9211 2658 9220
rect 2884 8566 2912 10066
rect 3160 9926 3188 10610
rect 3528 10554 3556 12174
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3436 10526 3556 10554
rect 3436 10062 3464 10526
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 1584 8288 1636 8294
rect 1306 8256 1362 8265
rect 1584 8230 1636 8236
rect 1306 8191 1362 8200
rect 1320 8090 1348 8191
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1596 7886 1624 8230
rect 2350 8188 2658 8197
rect 2350 8186 2356 8188
rect 2412 8186 2436 8188
rect 2492 8186 2516 8188
rect 2572 8186 2596 8188
rect 2652 8186 2658 8188
rect 2412 8134 2414 8186
rect 2594 8134 2596 8186
rect 2350 8132 2356 8134
rect 2412 8132 2436 8134
rect 2492 8132 2516 8134
rect 2572 8132 2596 8134
rect 2652 8132 2658 8134
rect 2350 8123 2658 8132
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1872 7546 1900 7822
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 2884 7478 2912 8502
rect 3436 8498 3464 9998
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2240 6866 2268 7414
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 3436 6798 3464 8434
rect 3528 8430 3556 10406
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3804 7342 3832 10134
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9722 3924 9862
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3896 8974 3924 9658
rect 3988 9110 4016 10406
rect 4080 10062 4108 11494
rect 4264 10674 4292 12038
rect 4356 11762 4384 12174
rect 4540 11762 4568 12582
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4896 12232 4948 12238
rect 5264 12232 5316 12238
rect 4948 12180 5120 12186
rect 4896 12174 5120 12180
rect 5264 12174 5316 12180
rect 4908 12158 5120 12174
rect 5092 12102 5120 12158
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 11694 4660 12038
rect 5092 11762 5120 12038
rect 5276 11898 5304 12174
rect 5368 11898 5396 12310
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4528 11552 4580 11558
rect 4448 11512 4528 11540
rect 4448 10674 4476 11512
rect 4528 11494 4580 11500
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4540 10674 4568 10950
rect 5276 10810 5304 11834
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4448 9926 4476 10610
rect 4540 10062 4568 10610
rect 5368 10470 5396 10610
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5460 10062 5488 13874
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5736 12918 5764 13262
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5552 12374 5580 12718
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5540 12232 5592 12238
rect 5644 12186 5672 12378
rect 5592 12180 5672 12186
rect 5540 12174 5672 12180
rect 5552 12158 5672 12174
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5552 10674 5580 11766
rect 5644 11694 5672 12038
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5736 10810 5764 12718
rect 5920 12374 5948 15506
rect 6472 15502 6500 17478
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 6012 14414 6040 14894
rect 6196 14482 6224 15370
rect 6288 14958 6316 15438
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6472 14550 6500 15438
rect 6564 14618 6592 18226
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6932 17202 6960 18022
rect 7116 17882 7144 18226
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7760 17338 7788 18226
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7852 17338 7880 17546
rect 8680 17542 8708 18226
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6656 16794 6684 17138
rect 6932 16794 6960 17138
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7760 16658 7788 17274
rect 8312 17202 8340 17478
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6748 15706 6776 16526
rect 8036 15706 8064 17138
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16794 8248 17070
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8220 16538 8248 16730
rect 8220 16510 8340 16538
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7932 15632 7984 15638
rect 7984 15580 8064 15586
rect 7932 15574 8064 15580
rect 7288 15564 7340 15570
rect 7944 15558 8064 15574
rect 7288 15506 7340 15512
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6748 15094 6776 15438
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6840 15042 6868 15302
rect 6932 15162 6960 15438
rect 7024 15162 7052 15438
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6460 14544 6512 14550
rect 6460 14486 6512 14492
rect 6184 14476 6236 14482
rect 6236 14436 6316 14464
rect 6184 14418 6236 14424
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6012 12850 6040 14350
rect 6104 12986 6132 14350
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 6104 12434 6132 12922
rect 6196 12442 6224 13806
rect 6288 12918 6316 14436
rect 6748 14414 6776 15030
rect 6840 15026 6960 15042
rect 6840 15020 6972 15026
rect 6840 15014 6920 15020
rect 6920 14962 6972 14968
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 14074 6408 14282
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 12714 6500 12786
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6012 12406 6132 12434
rect 6184 12436 6236 12442
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5828 11762 5856 12310
rect 6012 12238 6040 12406
rect 6184 12378 6236 12384
rect 6196 12322 6224 12378
rect 6104 12294 6224 12322
rect 6104 12238 6132 12294
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5816 11756 5868 11762
rect 6000 11756 6052 11762
rect 5868 11716 6000 11744
rect 5816 11698 5868 11704
rect 6000 11698 6052 11704
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5552 10266 5580 10474
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 5092 9874 5120 9998
rect 5092 9846 5212 9874
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3884 8968 3936 8974
rect 3936 8928 4016 8956
rect 3884 8910 3936 8916
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 7886 3924 8774
rect 3988 7886 4016 8928
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8498 4568 8774
rect 4816 8498 4844 8842
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4264 8022 4292 8434
rect 5184 8106 5212 9846
rect 5460 8498 5488 9998
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5552 8430 5580 10202
rect 5736 10062 5764 10746
rect 5828 10674 5856 11290
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 8974 5672 9862
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5644 8378 5672 8910
rect 5736 8634 5764 8978
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5724 8424 5776 8430
rect 5644 8372 5724 8378
rect 5644 8366 5776 8372
rect 5552 8242 5580 8366
rect 5644 8350 5764 8366
rect 5828 8362 5856 10610
rect 5920 10130 5948 10610
rect 6012 10538 6040 11698
rect 6104 11354 6132 12174
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6196 11898 6224 12106
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6472 11762 6500 12650
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6564 10606 6592 13738
rect 6748 12832 6776 14350
rect 6828 12844 6880 12850
rect 6748 12804 6828 12832
rect 6828 12786 6880 12792
rect 6932 10674 6960 14962
rect 7024 14958 7052 15098
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 13870 7144 14894
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12986 7052 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 10810 7144 12854
rect 7196 12232 7248 12238
rect 7300 12186 7328 15506
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 14482 7512 15302
rect 7576 15094 7604 15438
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7668 14958 7696 15438
rect 8036 15366 8064 15558
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7248 12180 7328 12186
rect 7196 12174 7328 12180
rect 7208 12158 7328 12174
rect 7208 11778 7236 12158
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11898 7328 12038
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7208 11750 7328 11778
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9722 5948 10066
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9722 6960 9998
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 5920 8498 5948 9658
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 8498 6684 8978
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 5552 8214 5672 8242
rect 5184 8078 5580 8106
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3896 6798 3924 7822
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 3804 5710 3832 6734
rect 3896 6458 3924 6734
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3988 5914 4016 6326
rect 4908 6322 4936 7346
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5460 6322 5488 6734
rect 5552 6322 5580 8078
rect 5644 6934 5672 8214
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5644 6798 5672 6870
rect 6564 6798 6592 8298
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 5552 5302 5580 6258
rect 5644 5370 5672 6258
rect 5828 5710 5856 6734
rect 6288 6390 6316 6734
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 6564 4690 6592 6734
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5778 6684 6054
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5234 6684 5510
rect 6840 5370 6868 8298
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6840 4554 6868 4966
rect 6932 4690 6960 9658
rect 7208 8974 7236 10474
rect 7300 10130 7328 11750
rect 7392 10810 7420 13194
rect 7576 12238 7604 14486
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7472 12232 7524 12238
rect 7564 12232 7616 12238
rect 7472 12174 7524 12180
rect 7562 12200 7564 12209
rect 7616 12200 7618 12209
rect 7484 12102 7512 12174
rect 7562 12135 7618 12144
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7392 9654 7420 10746
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 10266 7512 10542
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7104 8968 7156 8974
rect 7024 8928 7104 8956
rect 7024 8838 7052 8928
rect 7104 8910 7156 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7024 8498 7052 8774
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7024 7886 7052 8434
rect 7484 8294 7512 8978
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7116 6458 7144 7890
rect 7484 7886 7512 8230
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7576 7698 7604 10066
rect 7668 9722 7696 13806
rect 7760 11354 7788 14962
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7944 13530 7972 13874
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7840 12368 7892 12374
rect 7838 12336 7840 12345
rect 7932 12368 7984 12374
rect 7892 12336 7894 12345
rect 7932 12310 7984 12316
rect 7838 12271 7894 12280
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7760 10674 7788 11290
rect 7852 10674 7880 12038
rect 7944 11898 7972 12310
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7760 10538 7788 10610
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7760 9042 7788 10202
rect 8036 10062 8064 15302
rect 8128 15094 8156 15438
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 8312 13530 8340 16510
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13394 8432 14010
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8206 12336 8262 12345
rect 8206 12271 8262 12280
rect 8220 12238 8248 12271
rect 8208 12232 8260 12238
rect 8484 12232 8536 12238
rect 8208 12174 8260 12180
rect 8482 12200 8484 12209
rect 8536 12200 8538 12209
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7840 9036 7892 9042
rect 8036 9024 8064 9998
rect 7840 8978 7892 8984
rect 7944 8996 8064 9024
rect 7852 8498 7880 8978
rect 7944 8634 7972 8996
rect 8128 8974 8156 10474
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8036 8498 8064 8842
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7886 8064 8230
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7484 7670 7604 7698
rect 7484 7410 7512 7670
rect 8128 7546 8156 8910
rect 8220 8430 8248 12174
rect 8482 12135 8538 12144
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11762 8432 12038
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 9048 11014 9076 15370
rect 9324 14074 9352 18226
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9416 16810 9444 17138
rect 9508 16998 9536 17546
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9416 16782 9536 16810
rect 9508 16658 9536 16782
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 16114 9536 16594
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15162 9444 15982
rect 9508 15434 9536 16050
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9508 15162 9536 15370
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9416 14006 9444 15098
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9324 12986 9352 13194
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 8974 8340 10406
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9140 9586 9168 9930
rect 9324 9654 9352 11018
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9178 9260 9454
rect 9600 9450 9628 17138
rect 9692 16590 9720 18022
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10612 17202 10640 17478
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16114 9720 16526
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9968 15688 9996 17138
rect 10048 15700 10100 15706
rect 9968 15660 10048 15688
rect 9968 15366 9996 15660
rect 10048 15642 10100 15648
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 10704 15026 10732 18090
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10980 17338 11008 17546
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 9968 14822 9996 14962
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9968 13938 9996 14758
rect 10704 14414 10732 14962
rect 10980 14414 11008 16662
rect 11072 15570 11100 17546
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11348 15502 11376 15846
rect 11532 15502 11560 18022
rect 11900 17882 11928 18226
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11900 17202 11928 17818
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11348 15162 11376 15438
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11440 15162 11468 15302
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 14090 11008 14350
rect 10888 14062 11008 14090
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 9968 10674 9996 13874
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 10060 13258 10088 13806
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10796 13190 10824 13874
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12850 10824 13126
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10428 12481 10456 12786
rect 10414 12472 10470 12481
rect 10414 12407 10470 12416
rect 10796 12238 10824 12786
rect 10888 12782 10916 14062
rect 11164 13938 11192 14826
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14006 11376 14350
rect 11716 14074 11744 17138
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16794 11928 16934
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11992 15434 12020 15642
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 12176 15162 12204 15506
rect 12268 15434 12296 15846
rect 12544 15706 12572 18022
rect 13832 17066 13860 18022
rect 13924 17882 13952 18158
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13924 17338 13952 17818
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14292 17202 14320 17614
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 13096 15502 13124 16934
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13924 15706 13952 16050
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13648 15502 13676 15642
rect 14016 15638 14044 17138
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16182 14136 16934
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 14200 16114 14228 16390
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 13176 15496 13228 15502
rect 13544 15496 13596 15502
rect 13228 15444 13308 15450
rect 13176 15438 13308 15444
rect 13544 15438 13596 15444
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12636 14482 12664 15370
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11762 10640 12038
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10742 10732 11018
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 7546 8248 8366
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5234 7052 6054
rect 7116 5302 7144 6394
rect 7208 6254 7236 6734
rect 7484 6730 7512 7346
rect 8220 7002 8248 7482
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7484 6458 7512 6666
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7576 6458 7604 6598
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7484 6254 7512 6394
rect 7576 6322 7604 6394
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5710 7420 6054
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7116 5166 7144 5238
rect 8220 5234 8248 6802
rect 8956 6798 8984 7142
rect 9324 6866 9352 9114
rect 9876 9110 9904 9522
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 10152 8906 10180 9522
rect 10244 9178 10272 9522
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7478 9628 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9588 7336 9640 7342
rect 9508 7284 9588 7290
rect 9508 7278 9640 7284
rect 9508 7262 9628 7278
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8956 6322 8984 6734
rect 9140 6458 9168 6734
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 9140 5846 9168 6394
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 8128 5030 8156 5170
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6460 4548 6512 4554
rect 6460 4490 6512 4496
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 6472 4146 6500 4490
rect 6932 4146 6960 4626
rect 7944 4214 7972 4966
rect 8404 4622 8432 5510
rect 8392 4616 8444 4622
rect 8312 4564 8392 4570
rect 8312 4558 8444 4564
rect 8312 4542 8432 4558
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 8312 4078 8340 4542
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4214 8432 4422
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 9416 4146 9444 6190
rect 9508 5710 9536 7262
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 10244 5370 10272 7822
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 6866 10732 7346
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10336 5234 10364 5714
rect 10796 5250 10824 7686
rect 10888 6780 10916 10610
rect 10980 10266 11008 13874
rect 12820 13870 12848 14758
rect 12912 14618 12940 15302
rect 13096 15162 13124 15438
rect 13188 15422 13308 15438
rect 13280 15366 13308 15422
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13096 15026 13124 15098
rect 13280 15094 13308 15302
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13556 14958 13584 15438
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13740 15178 13768 15370
rect 13740 15150 13860 15178
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12912 14074 12940 14554
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13258 11836 13670
rect 13280 13546 13308 13874
rect 13832 13802 13860 15150
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 14004 13796 14056 13802
rect 14004 13738 14056 13744
rect 13280 13530 13400 13546
rect 13268 13524 13400 13530
rect 13320 13518 13400 13524
rect 13268 13466 13320 13472
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9586 11008 10066
rect 11072 9586 11100 11154
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 7546 11100 9522
rect 11256 9518 11284 10610
rect 11440 10130 11468 11630
rect 11808 10810 11836 12786
rect 12544 12442 12572 13194
rect 13280 12986 13308 13330
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13372 12850 13400 13518
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13832 12714 13860 13738
rect 14016 12850 14044 13738
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11992 11150 12020 11494
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 12084 11082 12112 11698
rect 12636 11354 12664 11698
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12728 11150 12756 11698
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11354 12848 11494
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12440 11008 12492 11014
rect 12820 10962 12848 11086
rect 12440 10950 12492 10956
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11256 7478 11284 9454
rect 11348 9450 11376 9862
rect 11440 9518 11468 10066
rect 11808 10062 11836 10746
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11808 9586 11836 9862
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11348 8498 11376 9386
rect 11440 8566 11468 9454
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11348 7954 11376 8434
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11440 7886 11468 8502
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11256 6866 11284 7414
rect 11440 7342 11468 7822
rect 11992 7818 12020 10406
rect 12452 9654 12480 10950
rect 12544 10934 12848 10962
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 9042 12480 9590
rect 12544 9382 12572 10934
rect 12912 10470 12940 11630
rect 13648 10810 13676 12650
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13740 10674 13768 11086
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 10968 6792 11020 6798
rect 10888 6752 10968 6780
rect 10968 6734 11020 6740
rect 10980 5574 11008 6734
rect 11256 6390 11284 6802
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5710 11376 6054
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10876 5296 10928 5302
rect 10704 5244 10876 5250
rect 10704 5238 10928 5244
rect 10704 5234 10916 5238
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10692 5228 10916 5234
rect 10744 5222 10916 5228
rect 10692 5170 10744 5176
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10152 4554 10180 4966
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 10980 4146 11008 5510
rect 11440 4622 11468 7278
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11808 6390 11836 6802
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 12452 6254 12480 7482
rect 12544 6798 12572 9318
rect 12728 9110 12756 9318
rect 13004 9178 13032 10406
rect 13832 10130 13860 12650
rect 14016 10470 14044 12786
rect 14108 12434 14136 15982
rect 14292 14090 14320 17138
rect 14936 16250 14964 17546
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15120 16114 15148 17002
rect 15672 16658 15700 17614
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14200 14062 14320 14090
rect 14384 14074 14412 14962
rect 14372 14068 14424 14074
rect 14200 12850 14228 14062
rect 14372 14010 14424 14016
rect 14476 13938 14504 15914
rect 14568 14482 14596 16050
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14752 15162 14780 15982
rect 15120 15314 15148 16050
rect 15672 15570 15700 16594
rect 16040 16114 16068 17478
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16592 16522 16620 16934
rect 16684 16658 16712 16934
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15120 15286 15240 15314
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15212 14958 15240 15286
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14292 13326 14320 13874
rect 14568 13802 14596 14418
rect 14936 13938 14964 14826
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14568 13326 14596 13738
rect 14660 13410 14688 13874
rect 14660 13382 14780 13410
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14108 12406 14228 12434
rect 14200 11694 14228 12406
rect 14476 12306 14504 13262
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14188 11688 14240 11694
rect 14188 11630 14240 11636
rect 14476 11082 14504 12242
rect 14568 12170 14596 12582
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12636 8634 12664 8910
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12820 8498 12848 8774
rect 13004 8498 13032 9114
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12636 8022 12664 8298
rect 13188 8090 13216 8366
rect 13464 8362 13492 8910
rect 13556 8906 13584 9386
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13924 8498 13952 9454
rect 14660 9450 14688 13194
rect 14752 12102 14780 13382
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11830 14780 12038
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14844 10810 14872 13874
rect 14936 13326 14964 13874
rect 15672 13394 15700 15506
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15856 15162 15884 15370
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15764 13326 15792 13670
rect 16040 13530 16068 14962
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 13938 16160 14894
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 14936 11694 14964 12718
rect 15028 12442 15056 12786
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15856 12238 15884 13330
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15580 11898 15608 12174
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 15948 11218 15976 12038
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15108 10600 15160 10606
rect 15028 10560 15108 10588
rect 15028 10130 15056 10560
rect 15108 10542 15160 10548
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15028 9518 15056 10066
rect 15120 9761 15148 10406
rect 15580 10062 15608 11086
rect 16132 10810 16160 11698
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16316 10606 16344 13738
rect 16776 12306 16804 17002
rect 16960 16454 16988 17070
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 17052 14618 17080 17138
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15745 17448 15846
rect 17406 15736 17462 15745
rect 17406 15671 17462 15680
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17236 14074 17264 15438
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17328 14958 17356 15302
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17236 13530 17264 13806
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17236 12918 17264 13466
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12345 16896 12582
rect 16854 12336 16910 12345
rect 16764 12300 16816 12306
rect 16854 12271 16910 12280
rect 16764 12242 16816 12248
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 10130 15884 10406
rect 16224 10266 16252 10542
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15106 9752 15162 9761
rect 15106 9687 15162 9696
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14016 8498 14044 9046
rect 15120 8974 15148 9687
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 13912 8492 13964 8498
rect 13832 8452 13912 8480
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5846 11744 6054
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11716 5710 11744 5782
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 12268 5166 12296 6190
rect 12544 6186 12572 6734
rect 12636 6662 12664 7958
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12820 6322 12848 6802
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5234 12388 5510
rect 12636 5370 12664 6258
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12728 5302 12756 6258
rect 12912 6118 12940 6598
rect 13556 6254 13584 6734
rect 13832 6458 13860 8452
rect 13912 8434 13964 8440
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14568 7478 14596 8774
rect 15580 7886 15608 9998
rect 16316 9042 16344 10542
rect 16408 9450 16436 12038
rect 16500 11354 16528 12038
rect 16776 11694 16804 12242
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16592 9654 16620 9930
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16868 9586 16896 12174
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16960 11082 16988 12038
rect 17328 11762 17356 14894
rect 17408 14408 17460 14414
rect 17406 14376 17408 14385
rect 17460 14376 17462 14385
rect 17406 14311 17462 14320
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17420 13705 17448 13874
rect 17406 13696 17462 13705
rect 17406 13631 17462 13640
rect 17406 13016 17462 13025
rect 17406 12951 17462 12960
rect 17420 12850 17448 12951
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17406 11656 17462 11665
rect 17406 11591 17408 11600
rect 17460 11591 17462 11600
rect 17408 11562 17460 11568
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 17406 10976 17462 10985
rect 17406 10911 17462 10920
rect 17420 10674 17448 10911
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17144 10305 17172 10610
rect 17130 10296 17186 10305
rect 17130 10231 17186 10240
rect 17406 9616 17462 9625
rect 16856 9580 16908 9586
rect 17406 9551 17408 9560
rect 16856 9522 16908 9528
rect 17460 9551 17462 9560
rect 17408 9522 17460 9528
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16408 8974 16436 9386
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16776 8838 16804 9454
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15580 7546 15608 7822
rect 15856 7546 15884 8774
rect 15948 7954 15976 8774
rect 16776 8430 16804 8774
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16776 8090 16804 8366
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7546 16804 7754
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 16868 7410 16896 9522
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15212 6914 15240 7278
rect 15120 6886 15240 6914
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12912 5098 12940 6054
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4826 12112 4966
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 13096 4690 13124 6190
rect 13832 4826 13860 6394
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14568 5914 14596 6326
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 15120 5710 15148 6886
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 14292 4622 14320 5646
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4282 11192 4490
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 14292 4146 14320 4558
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 16592 3602 16620 4150
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 17408 3528 17460 3534
rect 17406 3496 17408 3505
rect 17460 3496 17462 3505
rect 17406 3431 17462 3440
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
<< via2 >>
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 2356 17978 2412 17980
rect 2436 17978 2492 17980
rect 2516 17978 2572 17980
rect 2596 17978 2652 17980
rect 2356 17926 2402 17978
rect 2402 17926 2412 17978
rect 2436 17926 2466 17978
rect 2466 17926 2478 17978
rect 2478 17926 2492 17978
rect 2516 17926 2530 17978
rect 2530 17926 2542 17978
rect 2542 17926 2572 17978
rect 2596 17926 2606 17978
rect 2606 17926 2652 17978
rect 2356 17924 2412 17926
rect 2436 17924 2492 17926
rect 2516 17924 2572 17926
rect 2596 17924 2652 17926
rect 1306 17040 1362 17096
rect 846 14864 902 14920
rect 846 13096 902 13152
rect 2356 16890 2412 16892
rect 2436 16890 2492 16892
rect 2516 16890 2572 16892
rect 2596 16890 2652 16892
rect 2356 16838 2402 16890
rect 2402 16838 2412 16890
rect 2436 16838 2466 16890
rect 2466 16838 2478 16890
rect 2478 16838 2492 16890
rect 2516 16838 2530 16890
rect 2530 16838 2542 16890
rect 2542 16838 2572 16890
rect 2596 16838 2606 16890
rect 2606 16838 2652 16890
rect 2356 16836 2412 16838
rect 2436 16836 2492 16838
rect 2516 16836 2572 16838
rect 2596 16836 2652 16838
rect 2356 15802 2412 15804
rect 2436 15802 2492 15804
rect 2516 15802 2572 15804
rect 2596 15802 2652 15804
rect 2356 15750 2402 15802
rect 2402 15750 2412 15802
rect 2436 15750 2466 15802
rect 2466 15750 2478 15802
rect 2478 15750 2492 15802
rect 2516 15750 2530 15802
rect 2530 15750 2542 15802
rect 2542 15750 2572 15802
rect 2596 15750 2606 15802
rect 2606 15750 2652 15802
rect 2356 15748 2412 15750
rect 2436 15748 2492 15750
rect 2516 15748 2572 15750
rect 2596 15748 2652 15750
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 1398 10920 1454 10976
rect 2356 14714 2412 14716
rect 2436 14714 2492 14716
rect 2516 14714 2572 14716
rect 2596 14714 2652 14716
rect 2356 14662 2402 14714
rect 2402 14662 2412 14714
rect 2436 14662 2466 14714
rect 2466 14662 2478 14714
rect 2478 14662 2492 14714
rect 2516 14662 2530 14714
rect 2530 14662 2542 14714
rect 2542 14662 2572 14714
rect 2596 14662 2606 14714
rect 2606 14662 2652 14714
rect 2356 14660 2412 14662
rect 2436 14660 2492 14662
rect 2516 14660 2572 14662
rect 2596 14660 2652 14662
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 2356 13626 2412 13628
rect 2436 13626 2492 13628
rect 2516 13626 2572 13628
rect 2596 13626 2652 13628
rect 2356 13574 2402 13626
rect 2402 13574 2412 13626
rect 2436 13574 2466 13626
rect 2466 13574 2478 13626
rect 2478 13574 2492 13626
rect 2516 13574 2530 13626
rect 2530 13574 2542 13626
rect 2542 13574 2572 13626
rect 2596 13574 2606 13626
rect 2606 13574 2652 13626
rect 2356 13572 2412 13574
rect 2436 13572 2492 13574
rect 2516 13572 2572 13574
rect 2596 13572 2652 13574
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 2356 12538 2412 12540
rect 2436 12538 2492 12540
rect 2516 12538 2572 12540
rect 2596 12538 2652 12540
rect 2356 12486 2402 12538
rect 2402 12486 2412 12538
rect 2436 12486 2466 12538
rect 2466 12486 2478 12538
rect 2478 12486 2492 12538
rect 2516 12486 2530 12538
rect 2530 12486 2542 12538
rect 2542 12486 2572 12538
rect 2596 12486 2606 12538
rect 2606 12486 2652 12538
rect 2356 12484 2412 12486
rect 2436 12484 2492 12486
rect 2516 12484 2572 12486
rect 2596 12484 2652 12486
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 2356 11450 2412 11452
rect 2436 11450 2492 11452
rect 2516 11450 2572 11452
rect 2596 11450 2652 11452
rect 2356 11398 2402 11450
rect 2402 11398 2412 11450
rect 2436 11398 2466 11450
rect 2466 11398 2478 11450
rect 2478 11398 2492 11450
rect 2516 11398 2530 11450
rect 2530 11398 2542 11450
rect 2542 11398 2572 11450
rect 2596 11398 2606 11450
rect 2606 11398 2652 11450
rect 2356 11396 2412 11398
rect 2436 11396 2492 11398
rect 2516 11396 2572 11398
rect 2596 11396 2652 11398
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 2356 10362 2412 10364
rect 2436 10362 2492 10364
rect 2516 10362 2572 10364
rect 2596 10362 2652 10364
rect 2356 10310 2402 10362
rect 2402 10310 2412 10362
rect 2436 10310 2466 10362
rect 2466 10310 2478 10362
rect 2478 10310 2492 10362
rect 2516 10310 2530 10362
rect 2530 10310 2542 10362
rect 2542 10310 2572 10362
rect 2596 10310 2606 10362
rect 2606 10310 2652 10362
rect 2356 10308 2412 10310
rect 2436 10308 2492 10310
rect 2516 10308 2572 10310
rect 2596 10308 2652 10310
rect 2356 9274 2412 9276
rect 2436 9274 2492 9276
rect 2516 9274 2572 9276
rect 2596 9274 2652 9276
rect 2356 9222 2402 9274
rect 2402 9222 2412 9274
rect 2436 9222 2466 9274
rect 2466 9222 2478 9274
rect 2478 9222 2492 9274
rect 2516 9222 2530 9274
rect 2530 9222 2542 9274
rect 2542 9222 2572 9274
rect 2596 9222 2606 9274
rect 2606 9222 2652 9274
rect 2356 9220 2412 9222
rect 2436 9220 2492 9222
rect 2516 9220 2572 9222
rect 2596 9220 2652 9222
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 1306 8200 1362 8256
rect 2356 8186 2412 8188
rect 2436 8186 2492 8188
rect 2516 8186 2572 8188
rect 2596 8186 2652 8188
rect 2356 8134 2402 8186
rect 2402 8134 2412 8186
rect 2436 8134 2466 8186
rect 2466 8134 2478 8186
rect 2478 8134 2492 8186
rect 2516 8134 2530 8186
rect 2530 8134 2542 8186
rect 2542 8134 2572 8186
rect 2596 8134 2606 8186
rect 2606 8134 2652 8186
rect 2356 8132 2412 8134
rect 2436 8132 2492 8134
rect 2516 8132 2572 8134
rect 2596 8132 2652 8134
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 7562 12180 7564 12200
rect 7564 12180 7616 12200
rect 7616 12180 7618 12200
rect 7562 12144 7618 12180
rect 7838 12316 7840 12336
rect 7840 12316 7892 12336
rect 7892 12316 7894 12336
rect 7838 12280 7894 12316
rect 8206 12280 8262 12336
rect 8482 12180 8484 12200
rect 8484 12180 8536 12200
rect 8536 12180 8538 12200
rect 8482 12144 8538 12180
rect 10414 12416 10470 12472
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 17406 15680 17462 15736
rect 16854 12280 16910 12336
rect 15106 9696 15162 9752
rect 17406 14356 17408 14376
rect 17408 14356 17460 14376
rect 17460 14356 17462 14376
rect 17406 14320 17462 14356
rect 17406 13640 17462 13696
rect 17406 12960 17462 13016
rect 17406 11620 17462 11656
rect 17406 11600 17408 11620
rect 17408 11600 17460 11620
rect 17460 11600 17462 11620
rect 17406 10920 17462 10976
rect 17130 10240 17186 10296
rect 17406 9580 17462 9616
rect 17406 9560 17408 9580
rect 17408 9560 17460 9580
rect 17460 9560 17462 9580
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 17406 3476 17408 3496
rect 17408 3476 17460 3496
rect 17460 3476 17462 3496
rect 17406 3440 17462 3476
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
<< metal3 >>
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 3006 18463 3322 18464
rect 2346 17984 2662 17985
rect 2346 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2662 17984
rect 2346 17919 2662 17920
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 3006 17375 3322 17376
rect 0 17098 800 17128
rect 1301 17098 1367 17101
rect 0 17096 1367 17098
rect 0 17040 1306 17096
rect 1362 17040 1367 17096
rect 0 17038 1367 17040
rect 0 17008 800 17038
rect 1301 17035 1367 17038
rect 2346 16896 2662 16897
rect 2346 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2662 16896
rect 2346 16831 2662 16832
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 3006 16287 3322 16288
rect 2346 15808 2662 15809
rect 2346 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2662 15808
rect 2346 15743 2662 15744
rect 17401 15738 17467 15741
rect 18089 15738 18889 15768
rect 17401 15736 18889 15738
rect 17401 15680 17406 15736
rect 17462 15680 18889 15736
rect 17401 15678 18889 15680
rect 17401 15675 17467 15678
rect 18089 15648 18889 15678
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 3006 15199 3322 15200
rect 0 15058 800 15088
rect 0 14968 858 15058
rect 798 14925 858 14968
rect 798 14920 907 14925
rect 798 14864 846 14920
rect 902 14864 907 14920
rect 798 14862 907 14864
rect 841 14859 907 14862
rect 2346 14720 2662 14721
rect 2346 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2662 14720
rect 2346 14655 2662 14656
rect 17401 14378 17467 14381
rect 18089 14378 18889 14408
rect 17401 14376 18889 14378
rect 17401 14320 17406 14376
rect 17462 14320 18889 14376
rect 17401 14318 18889 14320
rect 17401 14315 17467 14318
rect 18089 14288 18889 14318
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 3006 14111 3322 14112
rect 17401 13698 17467 13701
rect 18089 13698 18889 13728
rect 17401 13696 18889 13698
rect 17401 13640 17406 13696
rect 17462 13640 18889 13696
rect 17401 13638 18889 13640
rect 17401 13635 17467 13638
rect 2346 13632 2662 13633
rect 2346 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2662 13632
rect 18089 13608 18889 13638
rect 2346 13567 2662 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 3006 13088 3322 13089
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 3006 13023 3322 13024
rect 17401 13018 17467 13021
rect 18089 13018 18889 13048
rect 17401 13016 18889 13018
rect 17401 12960 17406 13016
rect 17462 12960 18889 13016
rect 17401 12958 18889 12960
rect 0 12928 800 12958
rect 17401 12955 17467 12958
rect 18089 12928 18889 12958
rect 2346 12544 2662 12545
rect 2346 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2662 12544
rect 2346 12479 2662 12480
rect 10409 12474 10475 12477
rect 14958 12474 14964 12476
rect 10409 12472 14964 12474
rect 10409 12416 10414 12472
rect 10470 12416 14964 12472
rect 10409 12414 14964 12416
rect 10409 12411 10475 12414
rect 14958 12412 14964 12414
rect 15028 12412 15034 12476
rect 7833 12338 7899 12341
rect 8201 12338 8267 12341
rect 7833 12336 8267 12338
rect 7833 12280 7838 12336
rect 7894 12280 8206 12336
rect 8262 12280 8267 12336
rect 7833 12278 8267 12280
rect 7833 12275 7899 12278
rect 8201 12275 8267 12278
rect 16849 12338 16915 12341
rect 18089 12338 18889 12368
rect 16849 12336 18889 12338
rect 16849 12280 16854 12336
rect 16910 12280 18889 12336
rect 16849 12278 18889 12280
rect 16849 12275 16915 12278
rect 18089 12248 18889 12278
rect 7557 12202 7623 12205
rect 8477 12202 8543 12205
rect 7557 12200 8543 12202
rect 7557 12144 7562 12200
rect 7618 12144 8482 12200
rect 8538 12144 8543 12200
rect 7557 12142 8543 12144
rect 7557 12139 7623 12142
rect 8477 12139 8543 12142
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 3006 11935 3322 11936
rect 17401 11658 17467 11661
rect 18089 11658 18889 11688
rect 17401 11656 18889 11658
rect 17401 11600 17406 11656
rect 17462 11600 18889 11656
rect 17401 11598 18889 11600
rect 17401 11595 17467 11598
rect 18089 11568 18889 11598
rect 2346 11456 2662 11457
rect 2346 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2662 11456
rect 2346 11391 2662 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 17401 10978 17467 10981
rect 18089 10978 18889 11008
rect 17401 10976 18889 10978
rect 17401 10920 17406 10976
rect 17462 10920 18889 10976
rect 17401 10918 18889 10920
rect 17401 10915 17467 10918
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 18089 10888 18889 10918
rect 3006 10847 3322 10848
rect 2346 10368 2662 10369
rect 2346 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2662 10368
rect 2346 10303 2662 10304
rect 17125 10298 17191 10301
rect 18089 10298 18889 10328
rect 17125 10296 18889 10298
rect 17125 10240 17130 10296
rect 17186 10240 18889 10296
rect 17125 10238 18889 10240
rect 17125 10235 17191 10238
rect 18089 10208 18889 10238
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 3006 9759 3322 9760
rect 14958 9692 14964 9756
rect 15028 9754 15034 9756
rect 15101 9754 15167 9757
rect 15028 9752 15167 9754
rect 15028 9696 15106 9752
rect 15162 9696 15167 9752
rect 15028 9694 15167 9696
rect 15028 9692 15034 9694
rect 15101 9691 15167 9694
rect 17401 9618 17467 9621
rect 18089 9618 18889 9648
rect 17401 9616 18889 9618
rect 17401 9560 17406 9616
rect 17462 9560 18889 9616
rect 17401 9558 18889 9560
rect 17401 9555 17467 9558
rect 18089 9528 18889 9558
rect 2346 9280 2662 9281
rect 2346 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2662 9280
rect 2346 9215 2662 9216
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 2346 8192 2662 8193
rect 2346 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2662 8192
rect 2346 8127 2662 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 0 7488 800 7518
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 2346 4928 2662 4929
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 17401 3498 17467 3501
rect 18089 3498 18889 3528
rect 17401 3496 18889 3498
rect 17401 3440 17406 3496
rect 17462 3440 18889 3496
rect 17401 3438 18889 3440
rect 17401 3435 17467 3438
rect 18089 3408 18889 3438
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 2346 2687 2662 2688
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
<< via3 >>
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 2352 17980 2416 17984
rect 2352 17924 2356 17980
rect 2356 17924 2412 17980
rect 2412 17924 2416 17980
rect 2352 17920 2416 17924
rect 2432 17980 2496 17984
rect 2432 17924 2436 17980
rect 2436 17924 2492 17980
rect 2492 17924 2496 17980
rect 2432 17920 2496 17924
rect 2512 17980 2576 17984
rect 2512 17924 2516 17980
rect 2516 17924 2572 17980
rect 2572 17924 2576 17980
rect 2512 17920 2576 17924
rect 2592 17980 2656 17984
rect 2592 17924 2596 17980
rect 2596 17924 2652 17980
rect 2652 17924 2656 17980
rect 2592 17920 2656 17924
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 2352 16892 2416 16896
rect 2352 16836 2356 16892
rect 2356 16836 2412 16892
rect 2412 16836 2416 16892
rect 2352 16832 2416 16836
rect 2432 16892 2496 16896
rect 2432 16836 2436 16892
rect 2436 16836 2492 16892
rect 2492 16836 2496 16892
rect 2432 16832 2496 16836
rect 2512 16892 2576 16896
rect 2512 16836 2516 16892
rect 2516 16836 2572 16892
rect 2572 16836 2576 16892
rect 2512 16832 2576 16836
rect 2592 16892 2656 16896
rect 2592 16836 2596 16892
rect 2596 16836 2652 16892
rect 2652 16836 2656 16892
rect 2592 16832 2656 16836
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 2352 15804 2416 15808
rect 2352 15748 2356 15804
rect 2356 15748 2412 15804
rect 2412 15748 2416 15804
rect 2352 15744 2416 15748
rect 2432 15804 2496 15808
rect 2432 15748 2436 15804
rect 2436 15748 2492 15804
rect 2492 15748 2496 15804
rect 2432 15744 2496 15748
rect 2512 15804 2576 15808
rect 2512 15748 2516 15804
rect 2516 15748 2572 15804
rect 2572 15748 2576 15804
rect 2512 15744 2576 15748
rect 2592 15804 2656 15808
rect 2592 15748 2596 15804
rect 2596 15748 2652 15804
rect 2652 15748 2656 15804
rect 2592 15744 2656 15748
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 2352 14716 2416 14720
rect 2352 14660 2356 14716
rect 2356 14660 2412 14716
rect 2412 14660 2416 14716
rect 2352 14656 2416 14660
rect 2432 14716 2496 14720
rect 2432 14660 2436 14716
rect 2436 14660 2492 14716
rect 2492 14660 2496 14716
rect 2432 14656 2496 14660
rect 2512 14716 2576 14720
rect 2512 14660 2516 14716
rect 2516 14660 2572 14716
rect 2572 14660 2576 14716
rect 2512 14656 2576 14660
rect 2592 14716 2656 14720
rect 2592 14660 2596 14716
rect 2596 14660 2652 14716
rect 2652 14660 2656 14716
rect 2592 14656 2656 14660
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 2352 13628 2416 13632
rect 2352 13572 2356 13628
rect 2356 13572 2412 13628
rect 2412 13572 2416 13628
rect 2352 13568 2416 13572
rect 2432 13628 2496 13632
rect 2432 13572 2436 13628
rect 2436 13572 2492 13628
rect 2492 13572 2496 13628
rect 2432 13568 2496 13572
rect 2512 13628 2576 13632
rect 2512 13572 2516 13628
rect 2516 13572 2572 13628
rect 2572 13572 2576 13628
rect 2512 13568 2576 13572
rect 2592 13628 2656 13632
rect 2592 13572 2596 13628
rect 2596 13572 2652 13628
rect 2652 13572 2656 13628
rect 2592 13568 2656 13572
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 2352 12540 2416 12544
rect 2352 12484 2356 12540
rect 2356 12484 2412 12540
rect 2412 12484 2416 12540
rect 2352 12480 2416 12484
rect 2432 12540 2496 12544
rect 2432 12484 2436 12540
rect 2436 12484 2492 12540
rect 2492 12484 2496 12540
rect 2432 12480 2496 12484
rect 2512 12540 2576 12544
rect 2512 12484 2516 12540
rect 2516 12484 2572 12540
rect 2572 12484 2576 12540
rect 2512 12480 2576 12484
rect 2592 12540 2656 12544
rect 2592 12484 2596 12540
rect 2596 12484 2652 12540
rect 2652 12484 2656 12540
rect 2592 12480 2656 12484
rect 14964 12412 15028 12476
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 2352 11452 2416 11456
rect 2352 11396 2356 11452
rect 2356 11396 2412 11452
rect 2412 11396 2416 11452
rect 2352 11392 2416 11396
rect 2432 11452 2496 11456
rect 2432 11396 2436 11452
rect 2436 11396 2492 11452
rect 2492 11396 2496 11452
rect 2432 11392 2496 11396
rect 2512 11452 2576 11456
rect 2512 11396 2516 11452
rect 2516 11396 2572 11452
rect 2572 11396 2576 11452
rect 2512 11392 2576 11396
rect 2592 11452 2656 11456
rect 2592 11396 2596 11452
rect 2596 11396 2652 11452
rect 2652 11396 2656 11452
rect 2592 11392 2656 11396
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 2352 10364 2416 10368
rect 2352 10308 2356 10364
rect 2356 10308 2412 10364
rect 2412 10308 2416 10364
rect 2352 10304 2416 10308
rect 2432 10364 2496 10368
rect 2432 10308 2436 10364
rect 2436 10308 2492 10364
rect 2492 10308 2496 10364
rect 2432 10304 2496 10308
rect 2512 10364 2576 10368
rect 2512 10308 2516 10364
rect 2516 10308 2572 10364
rect 2572 10308 2576 10364
rect 2512 10304 2576 10308
rect 2592 10364 2656 10368
rect 2592 10308 2596 10364
rect 2596 10308 2652 10364
rect 2652 10308 2656 10364
rect 2592 10304 2656 10308
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 14964 9692 15028 9756
rect 2352 9276 2416 9280
rect 2352 9220 2356 9276
rect 2356 9220 2412 9276
rect 2412 9220 2416 9276
rect 2352 9216 2416 9220
rect 2432 9276 2496 9280
rect 2432 9220 2436 9276
rect 2436 9220 2492 9276
rect 2492 9220 2496 9276
rect 2432 9216 2496 9220
rect 2512 9276 2576 9280
rect 2512 9220 2516 9276
rect 2516 9220 2572 9276
rect 2572 9220 2576 9276
rect 2512 9216 2576 9220
rect 2592 9276 2656 9280
rect 2592 9220 2596 9276
rect 2596 9220 2652 9276
rect 2652 9220 2656 9276
rect 2592 9216 2656 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 2352 8188 2416 8192
rect 2352 8132 2356 8188
rect 2356 8132 2412 8188
rect 2412 8132 2416 8188
rect 2352 8128 2416 8132
rect 2432 8188 2496 8192
rect 2432 8132 2436 8188
rect 2436 8132 2492 8188
rect 2492 8132 2496 8188
rect 2432 8128 2496 8132
rect 2512 8188 2576 8192
rect 2512 8132 2516 8188
rect 2516 8132 2572 8188
rect 2572 8132 2576 8188
rect 2512 8128 2576 8132
rect 2592 8188 2656 8192
rect 2592 8132 2596 8188
rect 2596 8132 2652 8188
rect 2652 8132 2656 8188
rect 2592 8128 2656 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
<< metal4 >>
rect 2344 17984 2664 18544
rect 2344 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2664 17984
rect 2344 16896 2664 17920
rect 2344 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2664 16896
rect 2344 15808 2664 16832
rect 2344 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2664 15808
rect 2344 14720 2664 15744
rect 2344 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2664 14720
rect 2344 13632 2664 14656
rect 2344 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2664 13632
rect 2344 12544 2664 13568
rect 2344 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2664 12544
rect 2344 11456 2664 12480
rect 2344 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2664 11456
rect 2344 10368 2664 11392
rect 2344 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2664 10368
rect 2344 9280 2664 10304
rect 2344 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2664 9280
rect 2344 8192 2664 9216
rect 2344 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2664 8192
rect 2344 7104 2664 8128
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 3694 2664 3776
rect 2344 3458 2386 3694
rect 2622 3458 2664 3694
rect 2344 2752 2664 3458
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 2128 2664 2688
rect 3004 18528 3324 18544
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14176 3324 15200
rect 3004 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 14963 12476 15029 12477
rect 14963 12412 14964 12476
rect 15028 12412 15029 12476
rect 14963 12411 15029 12412
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 3004 8736 3324 9760
rect 14966 9757 15026 12411
rect 14963 9756 15029 9757
rect 14963 9692 14964 9756
rect 15028 9692 15029 9756
rect 14963 9691 15029 9692
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4354 3092 4384
rect 3156 4354 3172 4384
rect 3236 4354 3252 4384
rect 3316 4320 3324 4384
rect 3004 4118 3046 4320
rect 3282 4118 3324 4320
rect 3004 3296 3324 4118
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 2128 3324 2144
<< via4 >>
rect 2386 3458 2622 3694
rect 3046 4320 3076 4354
rect 3076 4320 3092 4354
rect 3092 4320 3156 4354
rect 3156 4320 3172 4354
rect 3172 4320 3236 4354
rect 3236 4320 3252 4354
rect 3252 4320 3282 4354
rect 3046 4118 3282 4320
<< metal5 >>
rect 1056 4354 17804 4396
rect 1056 4118 3046 4354
rect 3282 4118 17804 4354
rect 1056 4076 17804 4118
rect 1056 3694 17804 3736
rect 1056 3458 2386 3694
rect 2622 3458 17804 3694
rect 1056 3416 17804 3458
use sky130_fd_sc_hd__inv_2  _174_
timestamp -3599
transform -1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp -3599
transform -1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp -3599
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp -3599
transform -1 0 5888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp -3599
transform 1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp -3599
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp -3599
transform -1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp -3599
transform -1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp -3599
transform 1 0 11960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp -3599
transform -1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp -3599
transform -1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp -3599
transform -1 0 10672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _186_
timestamp -3599
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_4  _187_
timestamp -3599
transform 1 0 12420 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_4  _188_
timestamp -3599
transform -1 0 11408 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _189_
timestamp -3599
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp -3599
transform 1 0 2116 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _191_
timestamp -3599
transform 1 0 2024 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp -3599
transform 1 0 4140 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _193_
timestamp -3599
transform 1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _194_
timestamp -3599
transform 1 0 16008 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp -3599
transform 1 0 14444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _196_
timestamp -3599
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _197_
timestamp -3599
transform -1 0 13248 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand3b_4  _198_
timestamp -3599
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp -3599
transform 1 0 2116 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp -3599
transform 1 0 2208 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _202_
timestamp -3599
transform 1 0 4508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp -3599
transform 1 0 14720 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp -3599
transform 1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp -3599
transform 1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp -3599
transform 1 0 12144 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp -3599
transform -1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _208_
timestamp -3599
transform 1 0 11592 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp -3599
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _210_
timestamp -3599
transform -1 0 5428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _211_
timestamp -3599
transform 1 0 3864 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _212_
timestamp -3599
transform -1 0 5796 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _213_
timestamp -3599
transform 1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _214_
timestamp -3599
transform 1 0 3864 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _215_
timestamp -3599
transform -1 0 4048 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _216_
timestamp -3599
transform 1 0 4048 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _217_
timestamp -3599
transform 1 0 8096 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _218_
timestamp -3599
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _219_
timestamp -3599
transform 1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp -3599
transform -1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _221_
timestamp -3599
transform -1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _222_
timestamp -3599
transform -1 0 6072 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _223_
timestamp -3599
transform -1 0 14352 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _224_
timestamp -3599
transform -1 0 14076 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _225_
timestamp -3599
transform -1 0 13800 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _226_
timestamp -3599
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _227_
timestamp -3599
transform 1 0 12788 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _228_
timestamp -3599
transform 1 0 12052 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _229_
timestamp -3599
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _230_
timestamp -3599
transform -1 0 14076 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _231_
timestamp -3599
transform -1 0 14628 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _232_
timestamp -3599
transform -1 0 13616 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _233_
timestamp -3599
transform -1 0 13156 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_2  _234_
timestamp -3599
transform 1 0 12512 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _235_
timestamp -3599
transform -1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _236_
timestamp -3599
transform -1 0 8740 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _237_
timestamp -3599
transform -1 0 8464 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _238_
timestamp -3599
transform -1 0 8280 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _239_
timestamp -3599
transform -1 0 8004 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _240_
timestamp -3599
transform -1 0 7360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _241_
timestamp -3599
transform 1 0 6808 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp -3599
transform 1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _243_
timestamp -3599
transform 1 0 9568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _244_
timestamp -3599
transform 1 0 10028 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _245_
timestamp -3599
transform 1 0 12236 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _246_
timestamp -3599
transform -1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _247_
timestamp -3599
transform -1 0 11408 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _248_
timestamp -3599
transform -1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp -3599
transform -1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _250_
timestamp -3599
transform 1 0 12052 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _251_
timestamp -3599
transform 1 0 9292 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _252_
timestamp -3599
transform 1 0 10028 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _253_
timestamp -3599
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _254_
timestamp -3599
transform -1 0 9292 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _255_
timestamp -3599
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _256_
timestamp -3599
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_1  _257_
timestamp -3599
transform -1 0 9568 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _258_
timestamp -3599
transform -1 0 8740 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _259_
timestamp -3599
transform 1 0 7912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _260_
timestamp -3599
transform 1 0 6624 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _261_
timestamp -3599
transform -1 0 7728 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _262_
timestamp -3599
transform 1 0 5704 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _263_
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _264_
timestamp -3599
transform -1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _265_
timestamp -3599
transform 1 0 6072 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _266_
timestamp -3599
transform 1 0 5336 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _267_
timestamp -3599
transform 1 0 5152 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_1  _268_
timestamp -3599
transform 1 0 12696 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _269_
timestamp -3599
transform 1 0 12144 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _270_
timestamp -3599
transform 1 0 11500 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _271_
timestamp -3599
transform 1 0 12144 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _272_
timestamp -3599
transform -1 0 6164 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _273_
timestamp -3599
transform -1 0 5612 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _274_
timestamp -3599
transform -1 0 6992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _275_
timestamp -3599
transform -1 0 5980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _276_
timestamp -3599
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _277_
timestamp -3599
transform 1 0 7268 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp -3599
transform -1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _279_
timestamp -3599
transform -1 0 6256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _280_
timestamp -3599
transform -1 0 5704 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _281_
timestamp -3599
transform -1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _282_
timestamp -3599
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand4_1  _283_
timestamp -3599
transform 1 0 5060 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _284_
timestamp -3599
transform 1 0 7636 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _285_
timestamp -3599
transform 1 0 4324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _286_
timestamp -3599
transform 1 0 4048 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _287_
timestamp -3599
transform 1 0 4048 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _288_
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _289_
timestamp -3599
transform 1 0 3864 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _290_
timestamp -3599
transform -1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _291_
timestamp -3599
transform -1 0 9752 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _292_
timestamp -3599
transform -1 0 9844 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _293_
timestamp -3599
transform -1 0 9844 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _294_
timestamp -3599
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _295_
timestamp -3599
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _296_
timestamp -3599
transform 1 0 7912 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _297_
timestamp -3599
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _298_
timestamp -3599
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _299_
timestamp -3599
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp -3599
transform 1 0 7728 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _301_
timestamp -3599
transform 1 0 6992 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _302_
timestamp -3599
transform 1 0 7820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _303_
timestamp -3599
transform 1 0 6900 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _304_
timestamp -3599
transform 1 0 6256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _305_
timestamp -3599
transform 1 0 6532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _306_
timestamp -3599
transform 1 0 10948 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _307_
timestamp -3599
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _308_
timestamp -3599
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _309_
timestamp -3599
transform 1 0 14352 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _310_
timestamp -3599
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _311_
timestamp -3599
transform 1 0 15824 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp -3599
transform 1 0 14536 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _313_
timestamp -3599
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _314_
timestamp -3599
transform 1 0 15732 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp -3599
transform -1 0 14260 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _316_
timestamp -3599
transform -1 0 14444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _317_
timestamp -3599
transform 1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _318_
timestamp -3599
transform -1 0 13892 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _319_
timestamp -3599
transform 1 0 13800 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _320_
timestamp -3599
transform -1 0 15364 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp -3599
transform -1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _322_
timestamp -3599
transform -1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp -3599
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp -3599
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp -3599
transform -1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp -3599
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp -3599
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp -3599
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp -3599
transform 1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _330_
timestamp -3599
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp -3599
transform -1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp -3599
transform 1 0 12420 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp -3599
transform -1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp -3599
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp -3599
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp -3599
transform -1 0 5888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp -3599
transform -1 0 2852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp -3599
transform 1 0 4232 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp -3599
transform -1 0 3496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp -3599
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp -3599
transform 1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp -3599
transform 1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp -3599
transform 1 0 9936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp -3599
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp -3599
transform 1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp -3599
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp -3599
transform -1 0 3588 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _348_
timestamp -3599
transform -1 0 11132 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _349_
timestamp -3599
transform -1 0 3220 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _350_
timestamp -3599
transform -1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp -3599
transform 1 0 12144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _352_
timestamp -3599
transform 1 0 9292 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _353_
timestamp -3599
transform 1 0 13248 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _354_
timestamp -3599
transform 1 0 12052 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _355_
timestamp -3599
transform 1 0 9844 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _356_
timestamp -3599
transform 1 0 9016 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _357_
timestamp -3599
transform 1 0 7360 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _358_
timestamp -3599
transform -1 0 7268 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _359_
timestamp -3599
transform -1 0 4968 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _360_
timestamp -3599
transform 1 0 11500 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp -3599
transform 1 0 15548 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _362_
timestamp -3599
transform 1 0 15548 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp -3599
transform 1 0 14260 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp -3599
transform 1 0 3772 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _365_
timestamp -3599
transform 1 0 1564 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _366_
timestamp -3599
transform 1 0 3312 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp -3599
transform 1 0 1380 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp -3599
transform 1 0 15640 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _369_
timestamp -3599
transform -1 0 16008 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp -3599
transform 1 0 15640 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp -3599
transform 1 0 9016 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _372_
timestamp -3599
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _373_
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _374_
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _375_
timestamp -3599
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp -3599
transform 1 0 9200 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _377_
timestamp -3599
transform 1 0 7636 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _378_
timestamp -3599
transform 1 0 5704 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _379_
timestamp -3599
transform 1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _380_
timestamp -3599
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _381_
timestamp -3599
transform 1 0 10672 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _382_
timestamp -3599
transform 1 0 15916 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _383_
timestamp -3599
transform 1 0 15824 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _384_
timestamp -3599
transform 1 0 14628 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 8740 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -3599
transform -1 0 8188 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -3599
transform -1 0 7452 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -3599
transform 1 0 11776 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -3599
transform 1 0 11776 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp -3599
transform 1 0 5888 0 1 9792
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp -3599
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp -3599
transform 1 0 11776 0 -1 9792
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636964856
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636964856
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -3599
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636964856
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636964856
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -3599
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636964856
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636964856
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp -3599
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636964856
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636964856
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -3599
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636964856
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636964856
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp -3599
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636964856
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636964856
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -3599
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp -3599
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636964856
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636964856
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636964856
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636964856
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -3599
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -3599
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636964856
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636964856
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636964856
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636964856
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp -3599
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -3599
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp -3599
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp -3599
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636964856
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636964856
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636964856
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636964856
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636964856
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636964856
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp -3599
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636964856
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_153
timestamp -3599
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_161
timestamp -3599
transform 1 0 15916 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_60
timestamp -3599
transform 1 0 6624 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_91
timestamp 1636964856
transform 1 0 9476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp -3599
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -3599
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636964856
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636964856
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636964856
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636964856
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp -3599
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp -3599
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp -3599
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_41
timestamp -3599
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1636964856
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp -3599
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp -3599
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp -3599
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_118
timestamp -3599
transform 1 0 11960 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_144
timestamp 1636964856
transform 1 0 14352 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_156
timestamp 1636964856
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_168
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp -3599
transform 1 0 17296 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636964856
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636964856
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636964856
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636964856
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_66
timestamp -3599
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_83
timestamp 1636964856
transform 1 0 8740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp -3599
transform 1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp -3599
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_128
timestamp 1636964856
transform 1 0 12880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_140
timestamp 1636964856
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_152
timestamp 1636964856
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp -3599
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_169
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_177
timestamp -3599
transform 1 0 17388 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_33
timestamp 1636964856
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_45
timestamp -3599
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_49
timestamp -3599
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_55
timestamp 1636964856
transform 1 0 6164 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_67
timestamp 1636964856
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp -3599
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -3599
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp -3599
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_96
timestamp 1636964856
transform 1 0 9936 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_108
timestamp -3599
transform 1 0 11040 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_117
timestamp 1636964856
transform 1 0 11868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_129
timestamp -3599
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp -3599
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_148
timestamp 1636964856
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_160
timestamp 1636964856
transform 1 0 15824 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_172
timestamp -3599
transform 1 0 16928 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636964856
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_15
timestamp -3599
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp -3599
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp -3599
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_72
timestamp 1636964856
transform 1 0 7728 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_84
timestamp 1636964856
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_96
timestamp 1636964856
transform 1 0 9936 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp -3599
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_131
timestamp -3599
transform 1 0 13156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_155
timestamp 1636964856
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_177
timestamp -3599
transform 1 0 17388 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636964856
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_18
timestamp -3599
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp -3599
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_38
timestamp -3599
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp -3599
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_61
timestamp 1636964856
transform 1 0 6716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_73
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_88
timestamp 1636964856
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_100
timestamp -3599
transform 1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_106
timestamp 1636964856
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_118
timestamp -3599
transform 1 0 11960 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_128
timestamp 1636964856
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636964856
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636964856
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp -3599
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1636964856
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1636964856
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp -3599
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp -3599
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636964856
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp -3599
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp -3599
transform 1 0 8004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_79
timestamp -3599
transform 1 0 8372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_83
timestamp -3599
transform 1 0 8740 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636964856
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636964856
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp -3599
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_172
timestamp -3599
transform 1 0 16928 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_9
timestamp 1636964856
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp -3599
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -3599
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_35
timestamp 1636964856
transform 1 0 4324 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_47
timestamp 1636964856
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_59
timestamp -3599
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp -3599
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636964856
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_106
timestamp 1636964856
transform 1 0 10856 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_118
timestamp -3599
transform 1 0 11960 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_124
timestamp 1636964856
transform 1 0 12512 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp -3599
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636964856
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp -3599
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_26
timestamp -3599
transform 1 0 3496 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp -3599
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp -3599
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_65
timestamp -3599
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_78
timestamp 1636964856
transform 1 0 8280 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_90
timestamp 1636964856
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp -3599
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp -3599
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_118
timestamp -3599
transform 1 0 11960 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_147
timestamp 1636964856
transform 1 0 14628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp -3599
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp -3599
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_177
timestamp -3599
transform 1 0 17388 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636964856
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636964856
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -3599
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_35
timestamp 1636964856
transform 1 0 4324 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp -3599
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_54
timestamp -3599
transform 1 0 6072 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_68
timestamp -3599
transform 1 0 7360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -3599
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636964856
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636964856
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636964856
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_121
timestamp -3599
transform 1 0 12236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp -3599
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp -3599
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp -3599
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp -3599
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp -3599
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp -3599
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_171
timestamp -3599
transform 1 0 16836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp -3599
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636964856
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636964856
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636964856
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636964856
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp -3599
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp -3599
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_77
timestamp -3599
transform 1 0 8188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_102
timestamp -3599
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -3599
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp -3599
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_136
timestamp -3599
transform 1 0 13616 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_153
timestamp 1636964856
transform 1 0 15180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp -3599
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_172
timestamp -3599
transform 1 0 16928 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp -3599
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp -3599
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_37
timestamp -3599
transform 1 0 4508 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp -3599
transform 1 0 5060 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_51
timestamp -3599
transform 1 0 5796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp -3599
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636964856
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp -3599
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_105
timestamp -3599
transform 1 0 10764 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp -3599
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636964856
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp -3599
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp -3599
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_3
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_20
timestamp -3599
transform 1 0 2944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_28
timestamp -3599
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp -3599
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp -3599
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp -3599
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_75
timestamp -3599
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp -3599
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp -3599
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp -3599
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_121
timestamp -3599
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp -3599
transform 1 0 14352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_155
timestamp -3599
transform 1 0 15364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp -3599
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_6
timestamp 1636964856
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp -3599
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp -3599
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636964856
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636964856
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636964856
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636964856
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp -3599
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -3599
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp -3599
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_107
timestamp 1636964856
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_119
timestamp -3599
transform 1 0 12052 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_129
timestamp -3599
transform 1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp -3599
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636964856
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_153
timestamp -3599
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_157
timestamp -3599
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp -3599
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1636964856
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_40
timestamp -3599
transform 1 0 4784 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_48
timestamp -3599
transform 1 0 5520 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636964856
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp -3599
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_85
timestamp 1636964856
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_97
timestamp 1636964856
transform 1 0 10028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp -3599
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_132
timestamp 1636964856
transform 1 0 13248 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_144
timestamp -3599
transform 1 0 14352 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1636964856
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp -3599
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp -3599
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -3599
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_29
timestamp -3599
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_43
timestamp -3599
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_55
timestamp -3599
transform 1 0 6164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp -3599
transform 1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp -3599
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636964856
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp -3599
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp -3599
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_105
timestamp 1636964856
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_117
timestamp -3599
transform 1 0 11868 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_126
timestamp 1636964856
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp -3599
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp -3599
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636964856
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636964856
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp -3599
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp -3599
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_39
timestamp -3599
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_47
timestamp -3599
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp -3599
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1636964856
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1636964856
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_89
timestamp -3599
transform 1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp -3599
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp -3599
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_141
timestamp -3599
transform 1 0 14076 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_148
timestamp 1636964856
transform 1 0 14720 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp -3599
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp -3599
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_10
timestamp -3599
transform 1 0 2024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp -3599
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_38
timestamp -3599
transform 1 0 4600 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_46
timestamp -3599
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp -3599
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp -3599
transform 1 0 7820 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp -3599
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp -3599
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_106
timestamp -3599
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp -3599
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp -3599
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp -3599
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp -3599
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_151
timestamp -3599
transform 1 0 14996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_159
timestamp -3599
transform 1 0 15732 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp -3599
transform 1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp -3599
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp -3599
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp -3599
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_66
timestamp -3599
transform 1 0 7176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_70
timestamp -3599
transform 1 0 7544 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_87
timestamp -3599
transform 1 0 9108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_95
timestamp -3599
transform 1 0 9844 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp -3599
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -3599
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp -3599
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp -3599
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_129
timestamp -3599
transform 1 0 12972 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_135
timestamp -3599
transform 1 0 13524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_153
timestamp -3599
transform 1 0 15180 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp -3599
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp -3599
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp -3599
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp -3599
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1636964856
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp -3599
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_37
timestamp 1636964856
transform 1 0 4508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp -3599
transform 1 0 5612 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_61
timestamp 1636964856
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp -3599
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp -3599
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636964856
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_97
timestamp -3599
transform 1 0 10028 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_112
timestamp 1636964856
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 1636964856
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp -3599
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636964856
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636964856
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_165
timestamp -3599
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_173
timestamp -3599
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_6
timestamp -3599
transform 1 0 1656 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_21
timestamp 1636964856
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_33
timestamp -3599
transform 1 0 4140 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp -3599
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp -3599
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp -3599
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_72
timestamp 1636964856
transform 1 0 7728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_84
timestamp -3599
transform 1 0 8832 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_93
timestamp -3599
transform 1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp -3599
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp -3599
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_132
timestamp 1636964856
transform 1 0 13248 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_147
timestamp 1636964856
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_159
timestamp -3599
transform 1 0 15732 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp -3599
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp -3599
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp -3599
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp -3599
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp -3599
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_52
timestamp -3599
transform 1 0 5888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp -3599
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp -3599
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp -3599
transform 1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -3599
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_144
timestamp 1636964856
transform 1 0 14352 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp -3599
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_160
timestamp -3599
transform 1 0 15824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_177
timestamp -3599
transform 1 0 17388 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636964856
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp -3599
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_19
timestamp 1636964856
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_31
timestamp 1636964856
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_43
timestamp 1636964856
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp -3599
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636964856
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636964856
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_81
timestamp -3599
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp -3599
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1636964856
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp -3599
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp -3599
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636964856
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1636964856
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_137
timestamp -3599
transform 1 0 13708 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_145
timestamp -3599
transform 1 0 14444 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1636964856
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -3599
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp -3599
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636964856
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636964856
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -3599
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636964856
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636964856
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_53
timestamp -3599
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636964856
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp -3599
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp -3599
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp -3599
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_95
timestamp 1636964856
transform 1 0 9844 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_107
timestamp 1636964856
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_119
timestamp 1636964856
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp -3599
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -3599
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636964856
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_153
timestamp -3599
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_157
timestamp -3599
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp -3599
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_9
timestamp -3599
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_19
timestamp -3599
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_27
timestamp -3599
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_42
timestamp 1636964856
transform 1 0 4968 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp -3599
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_79
timestamp -3599
transform 1 0 8372 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp -3599
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_97
timestamp -3599
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_104
timestamp -3599
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_119
timestamp 1636964856
transform 1 0 12052 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_143
timestamp 1636964856
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_155
timestamp -3599
transform 1 0 15364 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_163
timestamp -3599
transform 1 0 16100 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp -3599
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp -3599
transform 1 0 7176 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp -3599
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_144
timestamp -3599
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_163
timestamp 1636964856
transform 1 0 16100 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_175
timestamp -3599
transform 1 0 17204 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp -3599
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1636964856
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_29
timestamp 1636964856
transform 1 0 3772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_41
timestamp -3599
transform 1 0 4876 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_49
timestamp -3599
transform 1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp -3599
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_63
timestamp -3599
transform 1 0 6900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp -3599
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_76
timestamp -3599
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_83
timestamp -3599
transform 1 0 8740 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp -3599
transform 1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_90
timestamp -3599
transform 1 0 9384 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_97
timestamp -3599
transform 1 0 10028 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp -3599
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -3599
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp -3599
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp -3599
transform 1 0 11960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp -3599
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp -3599
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_139
timestamp -3599
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_141
timestamp 1636964856
transform 1 0 14076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_153
timestamp 1636964856
transform 1 0 15180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp -3599
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp -3599
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp -3599
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3599
transform 1 0 11040 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input2
timestamp -3599
transform -1 0 17480 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3599
transform 1 0 13616 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3599
transform -1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -3599
transform -1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -3599
transform -1 0 10028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input7
timestamp -3599
transform -1 0 17480 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3599
transform -1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -3599
transform 1 0 17204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp -3599
transform 1 0 17204 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp -3599
transform -1 0 17204 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -3599
transform 1 0 5888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -3599
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp -3599
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp -3599
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -3599
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output17
timestamp -3599
transform -1 0 13248 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp -3599
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp -3599
transform -1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output20
timestamp -3599
transform 1 0 17204 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output21
timestamp -3599
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output22
timestamp -3599
transform 1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output23
timestamp -3599
transform -1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output24
timestamp -3599
transform -1 0 8096 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output25
timestamp -3599
transform -1 0 8740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output26
timestamp -3599
transform -1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output27
timestamp -3599
transform -1 0 9384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_30
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_31
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_32
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_33
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_34
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_35
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_36
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 17756 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_37
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_38
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 17756 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_39
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_40
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_41
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_42
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_43
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_44
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 17756 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_45
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 17756 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_46
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 17756 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_47
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_48
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 17756 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_49
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 17756 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_50
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_51
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_52
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 17756 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_53
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_54
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 17756 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_55
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_56
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 17756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_57
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_58
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 17756 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_59
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_67
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_70
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_73
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_76
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_91
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_100
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp -3599
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_103
timestamp -3599
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp -3599
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_106
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp -3599
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_109
timestamp -3599
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp -3599
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_112
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp -3599
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_115
timestamp -3599
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp -3599
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_118
timestamp -3599
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp -3599
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_121
timestamp -3599
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp -3599
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_124
timestamp -3599
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp -3599
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_127
timestamp -3599
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp -3599
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_130
timestamp -3599
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp -3599
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_133
timestamp -3599
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp -3599
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_136
timestamp -3599
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp -3599
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_139
timestamp -3599
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp -3599
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_142
timestamp -3599
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp -3599
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp -3599
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp -3599
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp -3599
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp -3599
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_150
timestamp -3599
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_151
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp -3599
transform 1 0 8832 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp -3599
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp -3599
transform 1 0 13984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_155
timestamp -3599
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
<< labels >>
flabel metal4 s 3004 2128 3324 18544 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4076 17804 4396 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2344 2128 2664 18544 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3416 17804 3736 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 10966 20233 11022 21033 0 FreeSans 224 90 0 0 addr[0]
port 2 nsew signal input
flabel metal3 s 18089 12928 18889 13048 0 FreeSans 480 0 0 0 addr[1]
port 3 nsew signal input
flabel metal2 s 13542 20233 13598 21033 0 FreeSans 224 90 0 0 addr[2]
port 4 nsew signal input
flabel metal2 s 12254 20233 12310 21033 0 FreeSans 224 90 0 0 addr[3]
port 5 nsew signal input
flabel metal3 s 18089 13608 18889 13728 0 FreeSans 480 0 0 0 addr[4]
port 6 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 clk
port 7 nsew signal input
flabel metal2 s 12898 20233 12954 21033 0 FreeSans 224 90 0 0 irq_timer
port 8 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 outa
port 9 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 outb
port 10 nsew signal output
flabel metal3 s 18089 15648 18889 15768 0 FreeSans 480 0 0 0 rdata[0]
port 11 nsew signal output
flabel metal3 s 18089 12248 18889 12368 0 FreeSans 480 0 0 0 rdata[1]
port 12 nsew signal output
flabel metal3 s 18089 11568 18889 11688 0 FreeSans 480 0 0 0 rdata[2]
port 13 nsew signal output
flabel metal2 s 11610 20233 11666 21033 0 FreeSans 224 90 0 0 rdata[3]
port 14 nsew signal output
flabel metal2 s 7746 20233 7802 21033 0 FreeSans 224 90 0 0 rdata[4]
port 15 nsew signal output
flabel metal2 s 8390 20233 8446 21033 0 FreeSans 224 90 0 0 rdata[5]
port 16 nsew signal output
flabel metal2 s 7102 20233 7158 21033 0 FreeSans 224 90 0 0 rdata[6]
port 17 nsew signal output
flabel metal2 s 9034 20233 9090 21033 0 FreeSans 224 90 0 0 rdata[7]
port 18 nsew signal output
flabel metal2 s 9678 20233 9734 21033 0 FreeSans 224 90 0 0 read_en
port 19 nsew signal input
flabel metal3 s 18089 3408 18889 3528 0 FreeSans 480 0 0 0 rst
port 20 nsew signal input
flabel metal3 s 18089 14288 18889 14408 0 FreeSans 480 0 0 0 wdata[0]
port 21 nsew signal input
flabel metal3 s 18089 10888 18889 11008 0 FreeSans 480 0 0 0 wdata[1]
port 22 nsew signal input
flabel metal3 s 18089 9528 18889 9648 0 FreeSans 480 0 0 0 wdata[2]
port 23 nsew signal input
flabel metal3 s 18089 10208 18889 10328 0 FreeSans 480 0 0 0 wdata[3]
port 24 nsew signal input
flabel metal2 s 5814 20233 5870 21033 0 FreeSans 224 90 0 0 wdata[4]
port 25 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 wdata[5]
port 26 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 wdata[6]
port 27 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 wdata[7]
port 28 nsew signal input
flabel metal2 s 10322 20233 10378 21033 0 FreeSans 224 90 0 0 write_en
port 29 nsew signal input
rlabel metal1 9430 18496 9430 18496 0 VGND
rlabel metal1 9430 17952 9430 17952 0 VPWR
rlabel metal2 9614 7582 9614 7582 0 _000_
rlabel metal1 13340 6358 13340 6358 0 _001_
rlabel metal1 12226 4794 12226 4794 0 _002_
rlabel metal2 10166 4760 10166 4760 0 _003_
rlabel metal1 9430 9622 9430 9622 0 _004_
rlabel metal1 7820 4182 7820 4182 0 _005_
rlabel metal1 6900 4522 6900 4522 0 _006_
rlabel metal1 4922 6222 4922 6222 0 _007_
rlabel metal1 3220 8398 3220 8398 0 _008_
rlabel metal2 3818 8738 3818 8738 0 _009_
rlabel metal2 14582 12376 14582 12376 0 _010_
rlabel metal2 16974 11560 16974 11560 0 _011_
rlabel metal2 10074 13532 10074 13532 0 _012_
rlabel metal1 4048 17306 4048 17306 0 _013_
rlabel metal1 2300 18054 2300 18054 0 _014_
rlabel metal2 2438 14110 2438 14110 0 _015_
rlabel metal1 3181 12138 3181 12138 0 _016_
rlabel metal2 9522 15266 9522 15266 0 _017_
rlabel metal1 2622 8568 2622 8568 0 _018_
rlabel metal1 2438 6834 2438 6834 0 _019_
rlabel metal1 13945 17578 13945 17578 0 _020_
rlabel metal2 10718 7106 10718 7106 0 _021_
rlabel metal2 14582 6120 14582 6120 0 _022_
rlabel metal1 13899 4522 13899 4522 0 _023_
rlabel metal1 11132 4250 11132 4250 0 _024_
rlabel metal2 10718 10880 10718 10880 0 _025_
rlabel metal2 8418 4318 8418 4318 0 _026_
rlabel metal2 6486 4318 6486 4318 0 _027_
rlabel metal2 4002 6120 4002 6120 0 _028_
rlabel metal2 12558 12818 12558 12818 0 _029_
rlabel metal1 16698 9622 16698 9622 0 _030_
rlabel metal2 16790 7650 16790 7650 0 _031_
rlabel metal1 16015 7446 16015 7446 0 _032_
rlabel metal1 5527 15402 5527 15402 0 _033_
rlabel metal2 2714 15640 2714 15640 0 _034_
rlabel metal1 4324 14246 4324 14246 0 _035_
rlabel metal1 3135 9962 3135 9962 0 _036_
rlabel metal1 16514 16966 16514 16966 0 _037_
rlabel metal2 15962 11628 15962 11628 0 _038_
rlabel metal1 9706 12954 9706 12954 0 _039_
rlabel metal2 4186 17476 4186 17476 0 _040_
rlabel metal1 1932 17306 1932 17306 0 _041_
rlabel metal1 1932 13498 1932 13498 0 _042_
rlabel metal1 1932 11866 1932 11866 0 _043_
rlabel metal2 9522 17272 9522 17272 0 _044_
rlabel metal2 7958 13702 7958 13702 0 _045_
rlabel via1 6021 17578 6021 17578 0 _046_
rlabel metal2 7866 17442 7866 17442 0 _047_
rlabel metal1 6624 16762 6624 16762 0 _048_
rlabel metal1 11270 17306 11270 17306 0 _049_
rlabel metal2 15870 15266 15870 15266 0 _050_
rlabel metal1 15952 13294 15952 13294 0 _051_
rlabel metal2 14950 16898 14950 16898 0 _052_
rlabel metal1 11224 15402 11224 15402 0 _053_
rlabel metal2 11822 13464 11822 13464 0 _054_
rlabel metal2 15870 10268 15870 10268 0 _055_
rlabel metal2 15962 8364 15962 8364 0 _056_
rlabel metal2 14582 8126 14582 8126 0 _057_
rlabel metal1 4462 15130 4462 15130 0 _058_
rlabel metal1 2116 15130 2116 15130 0 _059_
rlabel metal1 3772 13498 3772 13498 0 _060_
rlabel metal2 1702 10200 1702 10200 0 _061_
rlabel metal1 16330 16626 16330 16626 0 _062_
rlabel metal1 15042 11866 15042 11866 0 _063_
rlabel metal1 6762 9962 6762 9962 0 _064_
rlabel metal2 10626 11900 10626 11900 0 _065_
rlabel metal1 4968 12750 4968 12750 0 _066_
rlabel metal1 5750 12784 5750 12784 0 _067_
rlabel metal1 8004 8398 8004 8398 0 _068_
rlabel metal2 7498 12138 7498 12138 0 _069_
rlabel metal1 12650 9010 12650 9010 0 _070_
rlabel metal2 12834 11424 12834 11424 0 _071_
rlabel metal1 12972 11662 12972 11662 0 _072_
rlabel metal2 13110 16218 13110 16218 0 _073_
rlabel metal1 9522 17034 9522 17034 0 _074_
rlabel metal1 13156 15062 13156 15062 0 _075_
rlabel metal1 14766 13872 14766 13872 0 _076_
rlabel metal1 2438 17102 2438 17102 0 _077_
rlabel metal1 14582 14926 14582 14926 0 _078_
rlabel via1 2346 14909 2346 14909 0 _079_
rlabel metal1 11684 15130 11684 15130 0 _080_
rlabel metal2 12190 15334 12190 15334 0 _081_
rlabel metal1 4968 8466 4968 8466 0 _082_
rlabel metal2 4554 8636 4554 8636 0 _083_
rlabel metal2 5658 9418 5658 9418 0 _084_
rlabel metal1 5888 8602 5888 8602 0 _085_
rlabel metal2 4278 8228 4278 8228 0 _086_
rlabel metal1 4094 8500 4094 8500 0 _087_
rlabel metal1 5428 8874 5428 8874 0 _088_
rlabel metal1 7912 10234 7912 10234 0 _089_
rlabel metal1 6854 8908 6854 8908 0 _090_
rlabel metal2 7498 8058 7498 8058 0 _091_
rlabel metal1 6394 9010 6394 9010 0 _092_
rlabel metal2 12650 5814 12650 5814 0 _093_
rlabel metal2 9246 9316 9246 9316 0 _094_
rlabel metal1 13018 10608 13018 10608 0 _095_
rlabel metal1 13432 10778 13432 10778 0 _096_
rlabel metal1 13340 10642 13340 10642 0 _097_
rlabel metal1 13202 9146 13202 9146 0 _098_
rlabel metal2 12742 9214 12742 9214 0 _099_
rlabel metal2 13202 8228 13202 8228 0 _100_
rlabel metal2 12650 8772 12650 8772 0 _101_
rlabel metal1 13570 8534 13570 8534 0 _102_
rlabel metal1 13892 8398 13892 8398 0 _103_
rlabel metal2 13478 8636 13478 8636 0 _104_
rlabel metal1 12972 8806 12972 8806 0 _105_
rlabel metal1 12696 6086 12696 6086 0 _106_
rlabel metal2 10166 9214 10166 9214 0 _107_
rlabel metal1 7958 8908 7958 8908 0 _108_
rlabel metal1 7958 9010 7958 9010 0 _109_
rlabel metal2 8050 8058 8050 8058 0 _110_
rlabel metal1 7314 8908 7314 8908 0 _111_
rlabel metal2 9890 9316 9890 9316 0 _112_
rlabel metal2 7130 6528 7130 6528 0 _113_
rlabel metal1 9062 9418 9062 9418 0 _114_
rlabel metal1 9568 17170 9568 17170 0 _115_
rlabel metal2 12834 6562 12834 6562 0 _116_
rlabel metal1 11500 5678 11500 5678 0 _117_
rlabel metal1 11684 6086 11684 6086 0 _118_
rlabel metal2 12374 5372 12374 5372 0 _119_
rlabel metal2 10350 5474 10350 5474 0 _120_
rlabel metal1 10534 9554 10534 9554 0 _121_
rlabel metal2 8970 6970 8970 6970 0 _122_
rlabel metal1 9200 6834 9200 6834 0 _123_
rlabel metal1 9844 9486 9844 9486 0 _124_
rlabel metal2 8234 6018 8234 6018 0 _125_
rlabel metal1 6210 5746 6210 5746 0 _126_
rlabel metal1 6670 5678 6670 5678 0 _127_
rlabel metal2 6670 5372 6670 5372 0 _128_
rlabel metal1 5566 6800 5566 6800 0 _129_
rlabel metal1 5750 6698 5750 6698 0 _130_
rlabel metal2 5474 6528 5474 6528 0 _131_
rlabel metal1 12834 11866 12834 11866 0 _132_
rlabel metal2 12650 11526 12650 11526 0 _133_
rlabel metal1 12374 11696 12374 11696 0 _134_
rlabel metal1 8188 11730 8188 11730 0 _135_
rlabel metal2 5658 11866 5658 11866 0 _136_
rlabel metal2 5290 11322 5290 11322 0 _137_
rlabel metal1 4554 12240 4554 12240 0 _138_
rlabel metal1 5934 11866 5934 11866 0 _139_
rlabel metal2 7958 12104 7958 12104 0 _140_
rlabel metal1 4738 12172 4738 12172 0 _141_
rlabel metal1 4186 10608 4186 10608 0 _142_
rlabel metal1 7314 11662 7314 11662 0 _143_
rlabel metal1 5106 11696 5106 11696 0 _144_
rlabel metal2 8418 11900 8418 11900 0 _145_
rlabel metal1 7682 11764 7682 11764 0 _146_
rlabel metal1 4830 11594 4830 11594 0 _147_
rlabel metal1 4416 10642 4416 10642 0 _148_
rlabel metal2 4278 11356 4278 11356 0 _149_
rlabel metal1 4324 12614 4324 12614 0 _150_
rlabel metal2 4094 10778 4094 10778 0 _151_
rlabel metal1 9798 17034 9798 17034 0 _152_
rlabel metal2 15134 16558 15134 16558 0 _153_
rlabel metal2 14490 14926 14490 14926 0 _154_
rlabel metal1 6946 12886 6946 12886 0 _155_
rlabel metal2 7038 13124 7038 13124 0 _156_
rlabel metal2 6394 14178 6394 14178 0 _157_
rlabel metal1 6624 14586 6624 14586 0 _158_
rlabel metal1 7590 15402 7590 15402 0 _159_
rlabel metal1 7866 15674 7866 15674 0 _160_
rlabel metal2 6946 15300 6946 15300 0 _161_
rlabel metal1 6854 15674 6854 15674 0 _162_
rlabel metal2 10994 12070 10994 12070 0 _163_
rlabel metal1 11500 14042 11500 14042 0 _164_
rlabel metal1 14536 9418 14536 9418 0 _165_
rlabel metal1 15502 13498 15502 13498 0 _166_
rlabel metal1 14720 10778 14720 10778 0 _167_
rlabel metal1 15548 13906 15548 13906 0 _168_
rlabel metal2 14122 16558 14122 16558 0 _169_
rlabel metal2 14398 14518 14398 14518 0 _170_
rlabel metal1 14674 15130 14674 15130 0 _171_
rlabel metal1 13892 15674 13892 15674 0 _172_
rlabel metal1 14444 16218 14444 16218 0 _173_
rlabel metal1 10994 18258 10994 18258 0 addr[0]
rlabel metal2 17434 12903 17434 12903 0 addr[1]
rlabel metal2 13662 19295 13662 19295 0 addr[2]
rlabel metal2 12374 19295 12374 19295 0 addr[3]
rlabel metal2 17434 13787 17434 13787 0 addr[4]
rlabel metal3 1004 17068 1004 17068 0 clk
rlabel metal1 7774 9622 7774 9622 0 clknet_0_clk
rlabel metal1 7268 9690 7268 9690 0 clknet_2_0__leaf_clk
rlabel metal2 1426 13056 1426 13056 0 clknet_2_1__leaf_clk
rlabel metal1 13202 6222 13202 6222 0 clknet_2_2__leaf_clk
rlabel metal1 15916 12206 15916 12206 0 clknet_2_3__leaf_clk
rlabel metal1 13110 10472 13110 10472 0 cnt\[0\]
rlabel metal1 13018 6766 13018 6766 0 cnt\[1\]
rlabel metal1 14214 9486 14214 9486 0 cnt\[2\]
rlabel metal1 11638 11696 11638 11696 0 cnt\[3\]
rlabel metal1 7590 14994 7590 14994 0 cnt\[4\]
rlabel metal1 7774 15538 7774 15538 0 cnt\[5\]
rlabel metal1 6532 13838 6532 13838 0 cnt\[6\]
rlabel via1 5397 10642 5397 10642 0 cnt\[7\]
rlabel metal1 13662 11662 13662 11662 0 duty\[0\]
rlabel metal1 14858 11798 14858 11798 0 duty\[1\]
rlabel metal2 16514 11696 16514 11696 0 duty\[2\]
rlabel metal1 10672 12818 10672 12818 0 duty\[3\]
rlabel via2 7590 12189 7590 12189 0 duty\[4\]
rlabel metal1 2875 17510 2875 17510 0 duty\[5\]
rlabel metal1 4554 12886 4554 12886 0 duty\[6\]
rlabel via1 6486 12818 6486 12818 0 duty\[7\]
rlabel metal2 12742 5780 12742 5780 0 enable
rlabel metal2 13018 19363 13018 19363 0 irq_timer
rlabel metal1 12466 17544 12466 17544 0 irq_timer_next
rlabel metal1 13386 14926 13386 14926 0 net1
rlabel metal2 16422 10744 16422 10744 0 net10
rlabel metal2 15134 9333 15134 9333 0 net11
rlabel metal2 4554 17680 4554 17680 0 net12
rlabel metal1 2346 17170 2346 17170 0 net13
rlabel metal1 1610 13192 1610 13192 0 net14
rlabel metal1 2622 10778 2622 10778 0 net15
rlabel metal2 10718 16558 10718 16558 0 net16
rlabel metal2 13938 18020 13938 18020 0 net17
rlabel metal2 1610 8058 1610 8058 0 net18
rlabel metal1 1656 7514 1656 7514 0 net19
rlabel metal2 15088 10574 15088 10574 0 net2
rlabel metal1 16284 16082 16284 16082 0 net20
rlabel metal2 17250 13668 17250 13668 0 net21
rlabel metal1 17296 11730 17296 11730 0 net22
rlabel metal1 12006 17850 12006 17850 0 net23
rlabel metal2 7774 17782 7774 17782 0 net24
rlabel metal1 8556 17510 8556 17510 0 net25
rlabel via1 7130 18258 7130 18258 0 net26
rlabel metal1 9200 14042 9200 14042 0 net27
rlabel metal1 13662 17068 13662 17068 0 net3
rlabel metal1 13110 15674 13110 15674 0 net4
rlabel metal1 15778 15470 15778 15470 0 net5
rlabel metal1 9660 16558 9660 16558 0 net6
rlabel metal2 16606 3876 16606 3876 0 net7
rlabel metal1 17158 14586 17158 14586 0 net8
rlabel metal2 16146 11254 16146 11254 0 net9
rlabel metal1 1380 8058 1380 8058 0 outa
rlabel metal3 751 7548 751 7548 0 outb
rlabel metal2 13294 13702 13294 13702 0 period\[0\]
rlabel metal2 16238 10404 16238 10404 0 period\[1\]
rlabel metal2 16790 8228 16790 8228 0 period\[2\]
rlabel metal1 15548 8806 15548 8806 0 period\[3\]
rlabel metal1 7130 14994 7130 14994 0 period\[4\]
rlabel metal1 8096 15334 8096 15334 0 period\[5\]
rlabel metal1 5957 13906 5957 13906 0 period\[6\]
rlabel metal1 5252 10030 5252 10030 0 period\[7\]
rlabel metal2 17434 15793 17434 15793 0 rdata[0]
rlabel metal3 17488 12308 17488 12308 0 rdata[1]
rlabel via2 17434 11611 17434 11611 0 rdata[2]
rlabel metal2 11730 19363 11730 19363 0 rdata[3]
rlabel metal2 7866 19363 7866 19363 0 rdata[4]
rlabel metal2 8510 19363 8510 19363 0 rdata[5]
rlabel metal2 7222 19363 7222 19363 0 rdata[6]
rlabel metal2 9154 19363 9154 19363 0 rdata[7]
rlabel metal2 9982 19295 9982 19295 0 read_en
rlabel via2 17434 3485 17434 3485 0 rst
rlabel via2 17434 14365 17434 14365 0 wdata[0]
rlabel metal2 17434 10795 17434 10795 0 wdata[1]
rlabel via2 17434 9571 17434 9571 0 wdata[2]
rlabel metal2 17158 10455 17158 10455 0 wdata[3]
rlabel metal2 6118 19295 6118 19295 0 wdata[4]
rlabel metal3 751 15028 751 15028 0 wdata[5]
rlabel metal3 751 12988 751 12988 0 wdata[6]
rlabel metal3 1050 10948 1050 10948 0 wdata[7]
rlabel metal2 10534 19329 10534 19329 0 write_en
<< properties >>
string FIXED_BBOX 0 0 18889 21033
<< end >>
